* NGSPICE file created from egd_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

.subckt egd_top BitStream_buffer_input[0] BitStream_buffer_input[10] BitStream_buffer_input[11]
+ BitStream_buffer_input[12] BitStream_buffer_input[13] BitStream_buffer_input[14]
+ BitStream_buffer_input[15] BitStream_buffer_input[1] BitStream_buffer_input[2] BitStream_buffer_input[3]
+ BitStream_buffer_input[4] BitStream_buffer_input[5] BitStream_buffer_input[6] BitStream_buffer_input[7]
+ BitStream_buffer_input[8] BitStream_buffer_input[9] clk exp_golomb_decoding_output[0]
+ exp_golomb_decoding_output[1] exp_golomb_decoding_output[2] exp_golomb_decoding_output[3]
+ exp_golomb_decoding_output[4] exp_golomb_decoding_output[5] exp_golomb_decoding_output[6]
+ exp_golomb_decoding_output[7] exp_golomb_sel[0] exp_golomb_sel[1] half_fill_counter[0]
+ half_fill_counter[1] half_fill_counter[2] reset_counter[0] reset_counter[1] reset_counter[2]
+ reset_counter[3] reset_n vccd1 vssd1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3155_ _2688_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__buf_2
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3086_ BitStream_buffer.pc\[2\] _2604_ _2619_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__nor3_4
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3988_ BitStream_buffer.BS_buffer\[23\] _0351_ BitStream_buffer.BS_buffer\[24\] _0354_
+ _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__a221oi_1
X_5727_ _2351_ _2329_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5658_ net11 BitStream_buffer.BS_buffer\[123\] _2266_ vssd1 vssd1 vccd1 vccd1 _2291_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4609_ _3051_ _3034_ _3036_ _0521_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__a22o_1
X_5589_ _2243_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4960_ _1729_ _1733_ _1736_ _1738_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__and4_1
X_4891_ _3024_ _2848_ _1668_ _1669_ _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__o2111a_1
X_3911_ _0434_ _2744_ _0697_ _0698_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5512_ net1 BitStream_buffer.BS_buffer\[79\] _2156_ vssd1 vssd1 vccd1 vccd1 _2189_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3773_ _0551_ _0555_ _0559_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__and4_1
X_5443_ _2141_ _2127_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__and2_1
X_5374_ BitStream_buffer.pc_previous\[1\] BitStream_buffer.exp_golomb_len\[1\] vssd1
+ vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__or2_1
X_4325_ _2698_ _2670_ _0549_ _2675_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4256_ _2867_ _2829_ _1039_ _1040_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__o2111a_1
X_6014__112 clknet_1_0__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
X_4187_ _3027_ _3022_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__nor2_1
X_3207_ BitStream_buffer.BS_buffer\[94\] _2729_ BitStream_buffer.BS_buffer\[95\] _2732_
+ _2740_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__a221oi_1
X_3138_ _2641_ _2666_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__nand2_4
X_3069_ _2602_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5973__75 clknet_1_0__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__inv_2
X_6060__154 clknet_1_1__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__2584_ clknet_0__2584_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2584_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5090_ _2818_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__nand2_1
X_4110_ BitStream_buffer.BS_buffer\[79\] _2617_ BitStream_buffer.BS_buffer\[80\] _2624_
+ _0896_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4041_ _2835_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__nand2_1
X_4943_ _1691_ _1701_ _1722_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__nor3_1
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4874_ _2867_ _2779_ _1651_ _1652_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3825_ _2905_ _2916_ _2910_ _2920_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__o22ai_1
X_3756_ _0485_ _0545_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6109__39 clknet_1_0__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__inv_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3687_ _0400_ _2878_ BitStream_buffer.BS_buffer\[127\] _2876_ _0477_ vssd1 vssd1
+ vccd1 vccd1 _0478_ sky130_fd_sc_hd__a221oi_1
X_5426_ _2130_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
X_5357_ _2083_ _2079_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__and2_1
X_4308_ BitStream_buffer.BS_buffer\[22\] _0365_ BitStream_buffer.BS_buffer\[23\] _0369_
+ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__a221oi_1
X_5288_ net2 BitStream_buffer.BS_buffer\[37\] _2024_ vssd1 vssd1 vccd1 vccd1 _2036_
+ sky130_fd_sc_hd__mux2_1
X_4239_ _2733_ _2759_ _1022_ _1023_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3610_ _2904_ _0395_ _0401_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__nand3_1
X_4590_ BitStream_buffer.BS_buffer\[41\] _2929_ _2931_ BitStream_buffer.BS_buffer\[42\]
+ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__a22o_1
X_3541_ _3046_ _0332_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ net62 _0275_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[39\] sky130_fd_sc_hd__dfxtp_2
X_3472_ _2695_ _2965_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__and2_1
X_6191_ net153 _0206_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[85\] sky130_fd_sc_hd__dfxtp_1
X_5211_ _1976_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__clkbuf_1
X_5142_ _1914_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__nor2_1
X_5073_ _2748_ BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__nand2_1
X_4024_ _2765_ _2725_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4926_ _1702_ _1703_ _1704_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4857_ _2719_ _2816_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__nand2_1
X_3808_ _2856_ BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4788_ BitStream_buffer.BS_buffer\[1\] _2862_ _3039_ _2865_ _1568_ vssd1 vssd1 vccd1
+ vccd1 _1569_ sky130_fd_sc_hd__a221oi_1
Xclkbuf_0__2586_ _2586_ vssd1 vssd1 vccd1 vccd1 clknet_0__2586_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3739_ _0520_ _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5409_ net201 BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__nand2_1
X_6066__160 clknet_1_0__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5760_ _2329_ _2360_ BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1
+ vccd1 _2385_ sky130_fd_sc_hd__o21ai_1
X_5691_ _2315_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__inv_2
X_4711_ _1488_ _1490_ _1492_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4642_ _1422_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4573_ _0512_ _2852_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__or2_1
X_3524_ _3057_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__buf_2
X_6243_ net45 _0258_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[24\] sky130_fd_sc_hd__dfxtp_2
X_3455_ BitStream_buffer.BS_buffer\[48\] _2986_ _2988_ BitStream_buffer.BS_buffer\[49\]
+ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__a22o_1
X_6099__30 clknet_1_0__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__inv_2
X_3386_ _2919_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__buf_4
X_6174_ net136 _0189_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[102\] sky130_fd_sc_hd__dfxtp_1
X_5125_ BitStream_buffer.BS_buffer\[62\] _2985_ _2987_ BitStream_buffer.BS_buffer\[63\]
+ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__a22o_1
X_5056_ _2649_ BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4007_ _2625_ _2670_ _2631_ _2675_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__o22ai_1
X_5958_ _2560_ _2572_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__nand2_1
X_4909_ _0626_ _2954_ _0499_ _2958_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__o22ai_1
X_5889_ _2504_ _2475_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_5 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _2727_ _2741_ _2755_ _2773_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__and4_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _2639_ _2663_ _2684_ _2704_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5812_ _2322_ _2435_ _2348_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5743_ _2329_ _2360_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__nor2_1
X_5674_ _2121_ _2301_ _0675_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__a21oi_1
X_4625_ BitStream_buffer.BS_buffer\[37\] _0379_ BitStream_buffer.BS_buffer\[38\] _0383_
+ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4556_ _2870_ _2784_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__or2_1
X_3507_ _3040_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__buf_2
X_4487_ _0626_ _2941_ _0499_ _2945_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_40_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6226_ net188 _0241_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[50\] sky130_fd_sc_hd__dfxtp_4
X_3438_ BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__inv_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ net119 _0172_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[119\] sky130_fd_sc_hd__dfxtp_2
X_3369_ _2861_ _2874_ _2887_ _2902_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__and4_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _0604_ _2899_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__or2_1
X_5039_ BitStream_buffer.BS_buffer\[37\] _0336_ BitStream_buffer.BS_buffer\[38\] _0340_
+ _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[0] sky130_fd_sc_hd__buf_12
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 reset_counter[0] sky130_fd_sc_hd__buf_12
XFILLER_0_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6078__11 clknet_1_0__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__inv_2
XFILLER_0_37_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5979__81 clknet_1_0__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__inv_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4410_ _0388_ _0357_ _0654_ _0360_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5390_ _0405_ BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__nand2_1
X_4341_ _2761_ BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__nand2_1
X_4272_ _2953_ _2909_ _2956_ _2912_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o22ai_1
X_3223_ _2756_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__inv_2
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _2603_ _2687_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__nor2_2
X_3085_ _2618_ BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__nand2_4
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3987_ _0345_ _0357_ _0657_ _0360_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__o22ai_1
X_5726_ _2345_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__inv_4
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5657_ _2290_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4608_ _0523_ _3026_ _3053_ _3030_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__o22ai_1
X_5588_ _2242_ _2240_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__and2_1
X_4539_ _2756_ _2689_ _2725_ _2693_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__a221oi_1
X_6209_ net171 _0224_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[67\] sky130_fd_sc_hd__dfxtp_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4890_ _2858_ _0518_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__nand2_1
X_3910_ _0440_ _2753_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__or2_1
X_3841_ _0627_ _0628_ _0629_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3772_ BitStream_buffer.BS_buffer\[80\] _2689_ BitStream_buffer.BS_buffer\[81\] _2693_
+ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__a221oi_1
X_5511_ _2188_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5442_ net13 BitStream_buffer.BS_buffer\[57\] _2120_ vssd1 vssd1 vccd1 vccd1 _2141_
+ sky130_fd_sc_hd__mux2_1
X_5373_ _2094_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4324_ _0556_ _2646_ _1106_ _1107_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o2111a_1
X_4255_ _2894_ _2841_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__or2_1
X_4186_ _0968_ _0970_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__nand3b_1
X_3206_ _2733_ _2735_ _2737_ _2739_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__o22ai_1
X_3137_ BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__inv_2
X_3068_ _2600_ _2601_ BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5709_ _2333_ _1414_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6135__62 clknet_1_0__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__inv_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2583_ clknet_0__2583_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2583_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _2831_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__nand2_1
X_5991_ clknet_1_0__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__buf_1
X_4942_ _1712_ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4873_ _2790_ BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3824_ _0613_ _2909_ _0486_ _2912_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3755_ _0399_ BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3686_ _0476_ _2882_ _2880_ _2885_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5425_ _2129_ _2127_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5356_ net12 BitStream_buffer.BS_buffer\[26\] _2060_ vssd1 vssd1 vccd1 vccd1 _2083_
+ sky130_fd_sc_hd__mux2_1
X_5287_ _2035_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
X_4307_ _0657_ _0372_ _0534_ _0375_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__o22ai_1
X_4238_ _2715_ _2771_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__or2_1
X_4169_ BitStream_buffer.BS_buffer\[43\] _2924_ _2926_ BitStream_buffer.BS_buffer\[44\]
+ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3540_ _3052_ _3059_ _0324_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5210_ _1975_ _1973_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__and2_1
X_3471_ _3004_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__buf_2
X_6190_ net152 _0205_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[86\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6114__43 clknet_1_1__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__inv_2
X_5141_ _1915_ _1916_ _1917_ _1918_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5072_ _2745_ _2800_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__nand2_1
X_4023_ _2761_ _2721_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _0521_ _3040_ _3042_ BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1
+ _1705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4856_ _2811_ _2716_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3807_ _2845_ _2852_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__or2_1
X_4787_ _0730_ _2868_ _0604_ _2871_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_0__2585_ _2585_ vssd1 vssd1 vccd1 vccd1 clknet_0__2585_ sky130_fd_sc_hd__clkbuf_16
X_3738_ _0522_ _0524_ _0526_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3669_ _0459_ _2824_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__or2_1
X_5408_ _2116_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__inv_2
X_5339_ _2071_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5690_ _2314_ _0998_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__nand2_1
X_4710_ BitStream_buffer.BS_buffer\[70\] _3004_ BitStream_buffer.BS_buffer\[71\] _3007_
+ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4641_ BitStream_buffer.BS_buffer\[80\] _2678_ _2681_ BitStream_buffer.BS_buffer\[81\]
+ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4572_ _1342_ _1346_ _1350_ _1354_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__and4_1
X_3523_ _2943_ _3020_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__nand2_2
X_6242_ net44 _0257_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[25\] sky130_fd_sc_hd__dfxtp_2
X_3454_ _2987_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__buf_2
X_3385_ _2918_ _2907_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__nand2_2
X_6173_ net135 _0188_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[103\] sky130_fd_sc_hd__dfxtp_2
X_5124_ BitStream_buffer.BS_buffer\[68\] _2980_ _2982_ BitStream_buffer.BS_buffer\[69\]
+ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__a22o_1
X_5055_ _2725_ _2616_ _2706_ _2623_ _1832_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4006_ _2671_ _2646_ _0791_ _0792_ _0793_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _2569_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__inv_2
X_4908_ BitStream_buffer.BS_buffer\[56\] _2934_ BitStream_buffer.BS_buffer\[57\] _2937_
+ _1687_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__a221oi_1
X_5888_ _2504_ _2505_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4839_ _0398_ _0650_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_6 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ BitStream_buffer.BS_buffer\[78\] _2689_ BitStream_buffer.BS_buffer\[79\] _2693_
+ _2703_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5811_ _1310_ _2320_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5742_ _2366_ _1726_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5673_ _2118_ BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__nand2_1
X_4624_ _0739_ _0386_ _0613_ _0390_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__o22ai_1
X_4555_ _1327_ _1329_ _1333_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__and4_1
X_3506_ _3032_ _2648_ vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__nor2_2
X_4486_ _1266_ _1267_ _1268_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3437_ _2963_ _2967_ _2968_ _2970_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__o22ai_1
X_6225_ net187 _0240_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[51\] sky130_fd_sc_hd__dfxtp_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ net118 _0171_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[120\] sky130_fd_sc_hd__dfxtp_2
X_3368_ _2888_ _2890_ _2893_ _2897_ _2901_ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__o2111a_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _3018_ _2895_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__or2_1
X_3299_ _2831_ _2832_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__nand2_1
X_5038_ _0739_ _0343_ _0613_ _0346_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[1] sky130_fd_sc_hd__buf_12
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 reset_counter[1] sky130_fd_sc_hd__buf_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4340_ _0437_ _2744_ _1122_ _1123_ _1124_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o2111a_1
X_4271_ _1011_ _1026_ _1043_ _1056_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__and4_1
X_3222_ BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__clkbuf_4
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ _2647_ _2686_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__nand2_4
X_3084_ _2612_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__inv_2
X_3986_ BitStream_buffer.BS_buffer\[27\] _0337_ BitStream_buffer.BS_buffer\[28\] _0341_
+ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5725_ BitStream_buffer.BitStream_buffer_output\[5\] _2349_ vssd1 vssd1 vccd1 vccd1
+ _2350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5656_ _2289_ _2285_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4607_ _3063_ _3022_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__nor2_1
X_5587_ net2 BitStream_buffer.BS_buffer\[101\] _2230_ vssd1 vssd1 vccd1 vccd1 _2242_
+ sky130_fd_sc_hd__mux2_1
X_4538_ _0440_ _2697_ _2769_ _2702_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__o22ai_1
X_6069__2 clknet_1_1__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__inv_2
X_4469_ _2856_ _3039_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__nand2_1
X_6208_ net170 _0223_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[68\] sky130_fd_sc_hd__dfxtp_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3840_ BitStream_buffer.BS_buffer\[50\] _2986_ _2988_ BitStream_buffer.BS_buffer\[51\]
+ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3771_ _0560_ _2697_ _0419_ _2702_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_13_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5510_ _2187_ _2171_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ _2140_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
X_5372_ _2093_ _2079_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4323_ _0407_ _2661_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4254_ _2835_ BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__nand2_1
X_4185_ BitStream_buffer.BS_buffer\[65\] _3005_ BitStream_buffer.BS_buffer\[66\] _3008_
+ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__a221oi_1
X_3205_ _2738_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__buf_2
X_3136_ _2669_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__clkbuf_4
X_3067_ BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5708_ _2332_ _1518_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3969_ _2652_ _3011_ BitStream_buffer.BS_buffer\[66\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _0758_ sky130_fd_sc_hd__a2bb2o_1
X_5639_ net2 BitStream_buffer.BS_buffer\[117\] _2267_ vssd1 vssd1 vccd1 vccd1 _2278_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2582_ clknet_0__2582_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2582_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4941_ _1714_ _1716_ _1718_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__and4_1
X_4872_ _2786_ BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__nand2_1
X_3823_ BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3754_ _0498_ _0511_ _0544_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__nor3_1
XFILLER_0_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3685_ BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5424_ net4 BitStream_buffer.BS_buffer\[51\] _2121_ vssd1 vssd1 vccd1 vccd1 _2129_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5355_ _2082_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
X_5286_ _2033_ _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__and2_1
X_4306_ BitStream_buffer.BS_buffer\[26\] _0351_ BitStream_buffer.BS_buffer\[27\] _0354_
+ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__a221oi_1
X_4237_ _2765_ _2721_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4168_ _0739_ _2916_ _0613_ _2920_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__o22ai_1
X_4099_ _2914_ _0386_ _2917_ _0390_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__o22ai_1
X_3119_ _2642_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3470_ _2979_ _2699_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__nor2_2
XFILLER_0_51_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5140_ BitStream_buffer.BS_buffer\[23\] _0326_ _0328_ BitStream_buffer.BS_buffer\[22\]
+ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__a22o_1
X_5071_ _2832_ _2728_ _2838_ _2731_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__a221oi_1
X_4022_ _2769_ _2744_ _0807_ _0808_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__o2111a_1
X_4924_ _0363_ _3033_ _3035_ _0366_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4855_ _1625_ _1629_ _1632_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4786_ _3027_ _2848_ _1564_ _1565_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3806_ _0583_ _0587_ _0591_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__and4_1
X_3737_ _0527_ _0327_ _0329_ _0325_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2584_ _2584_ vssd1 vssd1 vccd1 vccd1 clknet_0__2584_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3668_ _2816_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
X_3599_ _0384_ _0386_ _0388_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__o22ai_1
X_5407_ _2618_ _0405_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__nand2_1
X_5338_ _2070_ _2055_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__and2_1
X_5269_ BitStream_buffer.buffer_index\[6\] _1946_ BitStream_buffer.buffer_index\[4\]
+ _1944_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__or4b_1
X_6027__124 clknet_1_0__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XFILLER_0_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4640_ _0560_ _2669_ _0419_ _2674_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4571_ _0727_ _2829_ _1351_ _1352_ _1353_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__o2111a_1
X_3522_ BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6241_ net43 _0256_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[26\] sky130_fd_sc_hd__dfxtp_2
X_3453_ _2654_ _2964_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__and2_2
X_6172_ net134 _0187_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[104\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3384_ _2648_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__inv_2
X_5123_ _2652_ _2973_ _2640_ _2976_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__o22ai_1
X_5054_ _2757_ _2629_ _0440_ _2636_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4005_ _0556_ _2661_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ _2570_ _2375_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5887_ _2448_ _2472_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__nor2_1
X_4907_ _2996_ _2940_ _2999_ _2944_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__o22ai_1
X_4838_ _1587_ _1597_ _1618_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__nor3_1
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4769_ _2870_ _2779_ _1547_ _1548_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5810_ _2432_ _2433_ _2393_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5741_ _2361_ _2328_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5672_ _2300_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4623_ BitStream_buffer.BS_buffer\[25\] _0365_ BitStream_buffer.BS_buffer\[26\] _0369_
+ _1405_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4554_ _0694_ _2759_ _1334_ _1335_ _1336_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__o2111a_1
X_3505_ BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4485_ BitStream_buffer.BS_buffer\[40\] _2929_ _2931_ BitStream_buffer.BS_buffer\[41\]
+ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6224_ net186 _0239_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[52\] sky130_fd_sc_hd__dfxtp_4
X_3436_ _2969_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__buf_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ net117 _0170_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[121\] sky130_fd_sc_hd__dfxtp_2
X_3367_ _2898_ _2900_ vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__or2_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _2891_ _0400_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__nand2_1
X_5037_ _1810_ _1815_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__nor2_1
X_3298_ BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5939_ _2505_ _2530_ _2504_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[2] sky130_fd_sc_hd__buf_12
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 reset_counter[2] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _1047_ _1049_ _1051_ _1055_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3221_ _2742_ _2744_ _2747_ _2750_ _2754_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__o2111a_1
X_3152_ _2685_ vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__inv_2
X_6084__16 clknet_1_0__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__inv_2
X_3083_ _2616_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3985_ _0388_ _0344_ _0654_ _0347_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__o22ai_1
X_5985__86 clknet_1_0__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__inv_2
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5724_ _2348_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5655_ net12 BitStream_buffer.BS_buffer\[122\] _2266_ vssd1 vssd1 vccd1 vccd1 _2289_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4606_ _1384_ _1386_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5586_ _2241_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4537_ _1318_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__nor2_1
X_4468_ _3018_ _2852_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__or2_1
X_6207_ net169 _0222_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[69\] sky130_fd_sc_hd__dfxtp_2
X_3419_ BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__inv_2
X_4399_ _0650_ _3034_ _3036_ _0770_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__a22o_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3770_ BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5440_ _2139_ _2127_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__and2_1
X_5371_ net1 BitStream_buffer.BS_buffer\[31\] _2060_ vssd1 vssd1 vccd1 vccd1 _2093_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ _2631_ _2656_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4253_ _2831_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3204_ _2700_ _2711_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__nand2_2
X_4184_ _2658_ _3011_ BitStream_buffer.BS_buffer\[68\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _0971_ sky130_fd_sc_hd__a2bb2o_1
X_3135_ _2668_ _2621_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__nand2_2
X_3066_ BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3968_ BitStream_buffer.BS_buffer\[59\] _2992_ BitStream_buffer.BS_buffer\[60\] _2995_
+ _0756_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__a221oi_1
X_5707_ _2331_ _1622_ vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__nand2_1
X_6071__4 clknet_1_1__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__inv_2
X_6021__119 clknet_1_1__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XFILLER_0_60_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3899_ BitStream_buffer.BS_buffer\[81\] _2689_ BitStream_buffer.BS_buffer\[82\] _2693_
+ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5638_ _2277_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5569_ _2228_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f__2581_ clknet_0__2581_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2581_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4940_ BitStream_buffer.BS_buffer\[40\] _0378_ BitStream_buffer.BS_buffer\[41\] _0382_
+ _1719_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4871_ _0601_ _2783_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3822_ _0563_ _0579_ _0596_ _0611_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__and4_1
X_3753_ _0530_ _0543_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3684_ BitStream_buffer.BS_buffer\[119\] _2863_ BitStream_buffer.BS_buffer\[120\]
+ _2866_ _0474_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__a221oi_1
X_5423_ _2128_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
X_5354_ _2081_ _2079_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__and2_1
X_4305_ _0654_ _0357_ _0531_ _0360_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__o22ai_1
X_5285_ _0404_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4236_ _2761_ _2736_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__nand2_1
X_4167_ _2956_ _2909_ _0847_ _2912_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3118_ BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__inv_2
X_4098_ BitStream_buffer.BS_buffer\[20\] _0365_ BitStream_buffer.BS_buffer\[21\] _0369_
+ _0885_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6004__103 clknet_1_0__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _2782_ _2734_ _0444_ _2738_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__o22ai_1
X_4021_ _2757_ _2753_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__or2_1
X_6050__145 clknet_1_0__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
X_4923_ _0370_ _3025_ _0373_ _3029_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4854_ _2721_ _2688_ _2714_ _2692_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4785_ _2858_ _3044_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__nand2_1
X_3805_ _2898_ _2829_ _0592_ _0593_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__o2111a_1
Xclkbuf_0__2583_ _2583_ vssd1 vssd1 vccd1 vccd1 clknet_0__2583_ sky130_fd_sc_hd__clkbuf_16
X_3736_ BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3667_ _2819_ BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__nand2_1
X_5406_ _2115_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
X_3598_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__buf_2
XFILLER_0_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5337_ net3 BitStream_buffer.BS_buffer\[20\] _2061_ vssd1 vssd1 vccd1 vccd1 _2070_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _2021_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
X_4219_ _0415_ _2646_ _1002_ _1003_ _1004_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__o2111a_1
X_5199_ net14 _0330_ _1950_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4570_ _0473_ _2841_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__or2_1
X_3521_ _3054_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6240_ net42 _0255_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[27\] sky130_fd_sc_hd__dfxtp_2
X_3452_ _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__clkbuf_4
X_3383_ BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__inv_2
X_6171_ net133 _0186_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[105\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5122_ _2658_ _2966_ _0411_ _2969_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__o22ai_1
X_5053_ _0672_ _1829_ _1831_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4004_ _2664_ _2656_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5955_ _2565_ _2569_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5886_ _2503_ _2415_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__nand2_2
X_4906_ _1682_ _1683_ _1684_ _1685_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__or4_1
X_4837_ _1608_ _1617_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4768_ _2790_ BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__nand2_1
X_4699_ _2963_ _2954_ _2968_ _2958_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3719_ BitStream_buffer.BS_buffer\[61\] _3005_ BitStream_buffer.BS_buffer\[62\] _3008_
+ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5740_ _2362_ _2364_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5671_ _2299_ _2285_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__and2_1
X_4622_ _0531_ _0372_ _0342_ _0375_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__o22ai_1
X_4553_ _0428_ _2771_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3504_ BitStream_buffer.BS_buffer\[4\] _3034_ _3036_ _3037_ vssd1 vssd1 vccd1 vccd1
+ _3038_ sky130_fd_sc_hd__a22o_1
X_4484_ BitStream_buffer.BS_buffer\[46\] _2924_ _2926_ BitStream_buffer.BS_buffer\[47\]
+ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__a22o_1
X_3435_ _2673_ _2965_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__nand2_2
X_6223_ net185 _0238_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[53\] sky130_fd_sc_hd__dfxtp_2
X_6056__151 clknet_1_1__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ net116 _0169_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[122\] sky130_fd_sc_hd__dfxtp_2
X_3366_ _2899_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__clkbuf_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _2830_ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__buf_2
X_5105_ _0770_ _2875_ _3051_ _2878_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__a221oi_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _1811_ _1812_ _1813_ _1814_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5938_ _2553_ _2375_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5869_ _2487_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.exp_golomb_len\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_31_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[3] sky130_fd_sc_hd__buf_12
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 reset_counter[3] sky130_fd_sc_hd__buf_12
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3220_ _2751_ _2753_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__or2_1
X_3151_ BitStream_buffer.pc\[2\] BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1
+ _2685_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3082_ _2603_ _2615_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3984_ _0766_ _0772_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5723_ _2329_ _2347_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5654_ _2288_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2589_ clknet_0__2589_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2589_
+ sky130_fd_sc_hd__clkbuf_16
X_4605_ BitStream_buffer.BS_buffer\[69\] _3005_ BitStream_buffer.BS_buffer\[70\] _3008_
+ _1387_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5585_ _2239_ _2240_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4536_ BitStream_buffer.BS_buffer\[79\] _2679_ _2682_ BitStream_buffer.BS_buffer\[80\]
+ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__a22o_1
X_4467_ _1238_ _1242_ _1246_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__and4_1
X_6206_ net168 _0221_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[70\] sky130_fd_sc_hd__dfxtp_2
X_4398_ _3056_ _3026_ _0648_ _3030_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__o22ai_1
X_3418_ _2951_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__buf_2
X_3349_ BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__inv_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ clknet_1_1__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__buf_1
X_5019_ BitStream_buffer.BS_buffer\[67\] _2980_ _2982_ BitStream_buffer.BS_buffer\[68\]
+ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5370_ _2092_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4321_ _2650_ BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4252_ _2839_ _2813_ _1035_ _1036_ _1037_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__o2111a_1
X_3203_ _2736_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ BitStream_buffer.BS_buffer\[61\] _2992_ BitStream_buffer.BS_buffer\[62\] _2995_
+ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__a221oi_1
X_3134_ _2667_ _2627_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__nor2_4
X_3065_ _2598_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _3009_ _2998_ _0632_ _3001_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5706_ _2330_ _1726_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3898_ _0686_ _2697_ _0560_ _2702_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5637_ _2276_ _2261_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5568_ _1945_ _1946_ BitStream_buffer.buffer_index\[4\] _1944_ vssd1 vssd1 vccd1
+ vccd1 _2228_ sky130_fd_sc_hd__or4b_2
XFILLER_0_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4519_ _0613_ _0386_ _0486_ _0390_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__o22ai_1
X_5499_ _2180_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__clkbuf_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__2580_ clknet_0__2580_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2580_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6126__54 clknet_1_1__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__inv_2
X_6141__68 clknet_1_1__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__inv_2
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4870_ _1639_ _1641_ _1645_ _1649_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__and4_1
X_3821_ _0600_ _0603_ _0606_ _0610_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3752_ _0533_ _0536_ _0539_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3683_ _0473_ _2869_ _2867_ _2872_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5422_ _2126_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__and2_1
X_5353_ net13 BitStream_buffer.BS_buffer\[25\] _2061_ vssd1 vssd1 vccd1 vccd1 _2081_
+ sky130_fd_sc_hd__mux2_1
X_4304_ _0387_ _0337_ BitStream_buffer.BS_buffer\[31\] _0341_ _1089_ vssd1 vssd1 vccd1
+ vccd1 _1090_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5284_ net3 BitStream_buffer.BS_buffer\[36\] _2024_ vssd1 vssd1 vccd1 vccd1 _2033_
+ sky130_fd_sc_hd__mux2_1
X_4235_ _2757_ _2744_ _1018_ _1019_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4166_ _0907_ _0922_ _0939_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3117_ _2650_ BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__nand2_1
X_4097_ _0355_ _0372_ _0358_ _0375_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4999_ _3063_ _2881_ _0640_ _2884_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _2749_ _2766_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__nand2_1
X_4922_ _0648_ _3021_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4853_ _2707_ _2696_ _0437_ _2701_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4784_ _2855_ _3037_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__nand2_1
X_3804_ _2827_ _2841_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__2582_ _2582_ vssd1 vssd1 vccd1 vccd1 clknet_0__2582_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3735_ _0525_ _3062_ _3060_ _0323_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5405_ _0405_ BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__nand2_1
X_3666_ _2815_ BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3597_ _2943_ _0338_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__nand2_2
X_5336_ _2069_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
X_6105__35 clknet_1_1__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__inv_2
X_5267_ _1986_ _1938_ _2020_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__a21o_1
X_6120__49 clknet_1_0__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__inv_2
X_4218_ _2625_ _2661_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__or2_1
X_5198_ _1967_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
X_4149_ _2835_ BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3520_ _2690_ _3020_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__nand2_2
X_3451_ _2979_ _2643_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__nor2_2
X_3382_ _2915_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__buf_2
X_6170_ net132 _0185_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[106\] sky130_fd_sc_hd__dfxtp_1
X_5121_ _1894_ _1896_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__nand3b_1
X_5052_ _1830_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4003_ _2650_ BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5954_ _2568_ _2415_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__nand2_1
X_5885_ _2497_ _2502_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__nand2_1
X_4905_ BitStream_buffer.BS_buffer\[44\] _2928_ _2930_ BitStream_buffer.BS_buffer\[45\]
+ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4836_ _1610_ _1612_ _1614_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4767_ _2786_ BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__nand2_1
X_4698_ BitStream_buffer.BS_buffer\[54\] _2934_ BitStream_buffer.BS_buffer\[55\] _2937_
+ _1479_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_43_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3718_ _0508_ _3011_ BitStream_buffer.BS_buffer\[64\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _0509_ sky130_fd_sc_hd__a2bb2o_1
X_3649_ _2762_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
X_5319_ net1 BitStream_buffer.BS_buffer\[47\] _2023_ vssd1 vssd1 vccd1 vccd1 _2057_
+ sky130_fd_sc_hd__mux2_1
X_6299_ net101 _0314_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_6033__130 clknet_1_1__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5670_ net1 BitStream_buffer.BS_buffer\[127\] _2266_ vssd1 vssd1 vccd1 vccd1 _2299_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4621_ _0380_ _0350_ _0387_ _0354_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__a221oi_1
X_4552_ _2765_ BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__nand2_1
X_3503_ BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__clkbuf_4
X_4483_ _2953_ _2916_ _2956_ _2920_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3434_ BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__inv_2
X_6222_ net184 _0237_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[54\] sky130_fd_sc_hd__dfxtp_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ net115 _0168_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[123\] sky130_fd_sc_hd__dfxtp_2
X_3365_ _2654_ _2847_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__nand2_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _3060_ _2881_ _3063_ _2884_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__o22ai_1
X_3296_ _2777_ _2699_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__nor2_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ BitStream_buffer.BS_buffer\[22\] _0326_ _0328_ BitStream_buffer.BS_buffer\[21\]
+ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5937_ _2550_ _2552_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5868_ _2608_ _2310_ _2327_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__or3_1
X_5799_ _2329_ _2360_ _1518_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__o21ai_1
X_4819_ BitStream_buffer.BS_buffer\[15\] _3033_ _3035_ _0363_ vssd1 vssd1 vccd1 vccd1
+ _1600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[4] sky130_fd_sc_hd__buf_12
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3150_ _2676_ _2683_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__nor2_1
X_3081_ _2614_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5722_ _2341_ _2345_ _2346_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__nand3_1
X_3983_ _0767_ _0768_ _0769_ _0771_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2588_ clknet_0__2588_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2588_
+ sky130_fd_sc_hd__clkbuf_16
X_5653_ _2287_ _2285_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4604_ _0556_ _3011_ BitStream_buffer.BS_buffer\[72\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _1387_ sky130_fd_sc_hd__a2bb2o_1
X_5584_ net19 vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4535_ _0419_ _2670_ _2694_ _2675_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4466_ _0601_ _2829_ _1247_ _1248_ _1249_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6205_ net167 _0220_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[71\] sky130_fd_sc_hd__dfxtp_2
X_4397_ _0514_ _3022_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nor2_1
X_3417_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3348_ _2881_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__buf_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _2812_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__buf_2
X_5018_ _2640_ _2973_ _0508_ _2976_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5990__91 clknet_1_1__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4320_ BitStream_buffer.BS_buffer\[81\] _2617_ BitStream_buffer.BS_buffer\[82\] _2624_
+ _1104_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__a221oi_1
X_4251_ _2782_ _2824_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__or2_1
X_3202_ BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4182_ _2640_ _2998_ _0508_ _3001_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__o22ai_1
X_3133_ _2666_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__inv_2
X_3064_ BitStream_buffer.BitStream_buffer_valid_n vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3966_ _0751_ _0752_ _0753_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5705_ _1830_ BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1 vccd1
+ _2330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5636_ net3 BitStream_buffer.BS_buffer\[116\] _2267_ vssd1 vssd1 vccd1 vccd1 _2276_
+ sky130_fd_sc_hd__mux2_1
X_3897_ BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5567_ _2227_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4518_ BitStream_buffer.BS_buffer\[24\] _0365_ BitStream_buffer.BS_buffer\[25\] _0369_
+ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__a221oi_1
X_5498_ _2179_ _2171_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__and2_1
X_4449_ _0568_ _2759_ _1230_ _1231_ _1232_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__o2111a_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3820_ _0481_ _2890_ _0607_ _0608_ _0609_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__o2111a_1
X_3751_ _0380_ _0379_ _0387_ _0383_ _0541_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3682_ BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5421_ _0404_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5352_ _2080_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4303_ _0663_ _0344_ _0540_ _0347_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5283_ _2032_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
X_4234_ _2707_ _2753_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4165_ _0943_ _0945_ _0947_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__and4_1
X_3116_ _2649_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__buf_2
X_4096_ BitStream_buffer.BS_buffer\[24\] _0351_ BitStream_buffer.BS_buffer\[25\] _0354_
+ _0883_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4998_ _3044_ _2862_ _0518_ _2865_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3949_ _0689_ _0705_ _0722_ _0737_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__and4_1
XFILLER_0_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5619_ _2263_ _2261_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4921_ _1696_ _1698_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__nand3b_1
X_4852_ _1630_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3803_ _2835_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__nand2_1
X_4783_ _0761_ _2851_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3734_ BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__inv_2
Xclkbuf_0__2581_ _2581_ vssd1 vssd1 vccd1 vccd1 clknet_0__2581_ sky130_fd_sc_hd__clkbuf_16
X_3665_ _2792_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5404_ _2611_ _2097_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc\[1\] sky130_fd_sc_hd__xor2_4
XFILLER_0_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3596_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__inv_2
X_5335_ _2068_ _2055_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__and2_1
X_5266_ _0673_ _2017_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _0556_ _2656_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__or2_1
X_5197_ _1966_ _1952_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__and2_1
X_4148_ _2831_ BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nand2_1
X_4079_ BitStream_buffer.BS_buffer\[64\] _3005_ BitStream_buffer.BS_buffer\[65\] _3008_
+ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3450_ BitStream_buffer.BS_buffer\[54\] _2981_ _2983_ BitStream_buffer.BS_buffer\[55\]
+ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3381_ _2659_ _2907_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__nand2_2
XFILLER_0_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ BitStream_buffer.BS_buffer\[54\] _2948_ BitStream_buffer.BS_buffer\[55\] _2951_
+ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__a221oi_1
X_5051_ BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1 vccd1 _1830_
+ sky130_fd_sc_hd__inv_2
X_4002_ BitStream_buffer.BS_buffer\[78\] _2617_ BitStream_buffer.BS_buffer\[79\] _2624_
+ _0789_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5953_ _2567_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5884_ _2498_ _2499_ _2349_ _2354_ _2501_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__o32a_1
XFILLER_0_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4904_ BitStream_buffer.BS_buffer\[50\] _2923_ _2925_ BitStream_buffer.BS_buffer\[51\]
+ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4835_ BitStream_buffer.BS_buffer\[39\] _0378_ BitStream_buffer.BS_buffer\[40\] _0382_
+ _1615_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4766_ _0473_ _2783_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3717_ BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4697_ _0858_ _2940_ _0750_ _2944_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3648_ _2765_ _2768_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__nand2_1
X_3579_ _2659_ _0338_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__nand2_2
X_5318_ _2056_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__clkbuf_1
X_6298_ net100 _0313_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_5249_ _2006_ _2007_ _0675_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096__27 clknet_1_0__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5997__97 clknet_1_1__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4620_ _0540_ _0357_ _0384_ _0360_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__o22ai_1
X_4551_ _2761_ BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3502_ _3035_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__buf_2
X_4482_ _0622_ _2909_ _0495_ _2912_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3433_ _2966_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__buf_2
X_6221_ net183 _0236_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[55\] sky130_fd_sc_hd__dfxtp_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ net114 _0167_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[124\] sky130_fd_sc_hd__dfxtp_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6017__115 clknet_1_0__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
X_3364_ BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__inv_2
X_5103_ _0518_ _2862_ _3037_ _2865_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__a221oi_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _2828_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__buf_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _0534_ _3061_ _0355_ _0322_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5936_ _2537_ _2538_ _2551_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__nand3_1
X_5867_ _2486_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.exp_golomb_len\[2\] sky130_fd_sc_hd__inv_2
X_6063__157 clknet_1_0__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XFILLER_0_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5798_ _2370_ _2390_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__nand2_1
X_4818_ _0373_ _3025_ _0646_ _3029_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__o22ai_1
X_4749_ _2706_ _2688_ _2721_ _2692_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__a221oi_1
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[5] sky130_fd_sc_hd__buf_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3080_ BitStream_buffer.pc\[2\] _2604_ _2613_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _0770_ _0327_ _0329_ _0650_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__a22o_1
X_5721_ BitStream_buffer.BitStream_buffer_output\[15\] BitStream_buffer.BitStream_buffer_valid_n
+ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5652_ net13 BitStream_buffer.BS_buffer\[121\] _2267_ vssd1 vssd1 vccd1 vccd1 _2287_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__2587_ clknet_0__2587_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2587_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4603_ BitStream_buffer.BS_buffer\[65\] _2992_ BitStream_buffer.BS_buffer\[66\] _2995_
+ _1385_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__a221oi_1
X_5583_ net3 _2820_ _2230_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4534_ _2625_ _2646_ _1314_ _1315_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__o2111a_1
X_4465_ _2867_ _2841_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__or2_1
X_3416_ _2628_ _2907_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__and2_1
X_4396_ _1176_ _1178_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__nand3b_1
X_6204_ net166 _0219_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[72\] sky130_fd_sc_hd__dfxtp_2
X_3347_ _2695_ _2847_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__nand2_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3278_ _2680_ _2778_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__nand2_2
X_5017_ _0411_ _2966_ _2652_ _2969_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5976__78 clknet_1_0__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__inv_2
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5919_ _2534_ _2535_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__nand2_1
XFILLER_0_8_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _2819_ _2788_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__nand2_1
X_4181_ _0964_ _0965_ _0966_ _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__or4_1
X_3201_ _2734_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__buf_2
X_3132_ BitStream_buffer.pc\[3\] _2665_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3965_ BitStream_buffer.BS_buffer\[51\] _2986_ _2988_ BitStream_buffer.BS_buffer\[52\]
+ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5704_ _2328_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__inv_6
X_3896_ _0683_ _0684_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5635_ _2275_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5566_ _2226_ _2216_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4517_ _0342_ _0372_ _0345_ _0375_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__o22ai_1
X_5497_ net12 BitStream_buffer.BS_buffer\[74\] _2156_ vssd1 vssd1 vccd1 vccd1 _2179_
+ sky130_fd_sc_hd__mux2_1
X_4448_ _2733_ _2771_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__or2_1
X_4379_ BitStream_buffer.BS_buffer\[45\] _2924_ _2926_ BitStream_buffer.BS_buffer\[46\]
+ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__a22o_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3750_ _0540_ _0386_ _0384_ _0390_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3681_ _2883_ _2849_ _0469_ _0470_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5420_ net5 BitStream_buffer.BS_buffer\[50\] _2121_ vssd1 vssd1 vccd1 vccd1 _2126_
+ sky130_fd_sc_hd__mux2_1
X_5351_ _2078_ _2079_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5282_ _2031_ _1973_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4302_ _1082_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__nor2_1
X_4233_ _2749_ _2762_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__nand2_1
X_4164_ _2867_ _2890_ _0948_ _0949_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__o2111a_1
X_4095_ _0342_ _0357_ _0345_ _0360_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3115_ _2603_ _2648_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__nor2_2
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _0512_ _2868_ _3018_ _2871_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3948_ _0726_ _0729_ _0732_ _0736_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3879_ _0399_ _3039_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__nand2_1
X_5618_ net1 BitStream_buffer.BS_buffer\[111\] _2229_ vssd1 vssd1 vccd1 vccd1 _2263_
+ sky130_fd_sc_hd__mux2_1
X_5549_ net12 _2721_ _2192_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ BitStream_buffer.BS_buffer\[72\] _3004_ BitStream_buffer.BS_buffer\[73\] _3007_
+ _1699_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4851_ BitStream_buffer.BS_buffer\[82\] _2678_ _2681_ BitStream_buffer.BS_buffer\[83\]
+ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3802_ _2831_ _2836_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__nand2_1
X_4782_ _1550_ _1554_ _1558_ _1562_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2580_ _2580_ vssd1 vssd1 vccd1 vccd1 clknet_0__2580_ sky130_fd_sc_hd__clkbuf_16
X_3733_ _0523_ _3055_ _3053_ _3058_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_55_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3664_ _0450_ _2797_ _0451_ _0452_ _0454_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__o2111a_1
X_5403_ _2114_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3595_ BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5334_ net4 BitStream_buffer.BS_buffer\[19\] _2061_ vssd1 vssd1 vccd1 vccd1 _2068_
+ sky130_fd_sc_hd__mux2_1
X_5265_ _2019_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__clkbuf_1
X_5196_ net15 BitStream_buffer.BS_buffer\[7\] _1950_ vssd1 vssd1 vccd1 vccd1 _1966_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4216_ _2650_ BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__nand2_1
X_4147_ _0445_ _2813_ _0931_ _0932_ _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__o2111a_1
X_4078_ _0411_ _3011_ BitStream_buffer.BS_buffer\[67\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _0866_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3380_ BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__inv_2
X_5050_ _1785_ _1827_ _1828_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__nand3_1
X_4001_ _2694_ _2630_ _2698_ _2637_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__o22ai_1
X_6110__40 clknet_1_0__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__inv_2
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5952_ _2566_ _2381_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4903_ _2939_ _2915_ _2942_ _2919_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5883_ BitStream_buffer.BitStream_buffer_output\[11\] _2500_ vssd1 vssd1 vccd1 vccd1
+ _2501_ sky130_fd_sc_hd__xor2_1
X_4834_ _2956_ _0385_ _0847_ _0389_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__o22ai_1
X_4765_ _1535_ _1537_ _1541_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__and4_1
X_3716_ BitStream_buffer.BS_buffer\[57\] _2992_ BitStream_buffer.BS_buffer\[58\] _2995_
+ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4696_ _1474_ _1475_ _1476_ _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__or4_1
X_3647_ _2761_ _2756_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__nand2_1
X_3578_ BitStream_buffer.BS_buffer\[19\] vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5317_ _2054_ _2055_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__and2_1
X_6297_ net99 _0312_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_5248_ _2001_ net29 vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__nand2_1
X_5179_ _1954_ _1952_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6040__136 clknet_1_1__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4550_ _0423_ _2744_ _1330_ _1331_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3501_ _2668_ _3020_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__and2_2
X_4481_ _1219_ _1234_ _1251_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__and4_1
X_3432_ _2668_ _2965_ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__nand2_2
X_6220_ net182 _0235_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[56\] sky130_fd_sc_hd__dfxtp_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ net113 _0166_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[125\] sky130_fd_sc_hd__dfxtp_2
X_3363_ _2894_ _2896_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__or2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5102_ _0638_ _2868_ _0512_ _2871_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__o22ai_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _2690_ _2778_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__nand2_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _0531_ _3054_ _0342_ _3057_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6074__7 clknet_1_0__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__inv_2
X_5935_ _2549_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5866_ _2608_ _2310_ _2345_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__or3_1
X_4817_ _0525_ _3021_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__nor2_1
X_5797_ _2308_ net18 _2309_ _2606_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _0437_ _2696_ _2757_ _2701_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__o22ai_1
X_4679_ _2855_ _0518_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[6] sky130_fd_sc_hd__buf_12
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__clkbuf_4
X_5720_ _2343_ _2318_ _2344_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2586_ clknet_0__2586_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2586_
+ sky130_fd_sc_hd__clkbuf_16
X_5651_ _2286_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4602_ _2671_ _2998_ _2658_ _3001_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__o22ai_1
X_5582_ _2238_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4533_ _2698_ _2661_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _2835_ BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__nand2_1
X_6203_ net165 _0218_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[73\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3415_ _2948_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__buf_2
X_4395_ BitStream_buffer.BS_buffer\[67\] _3005_ BitStream_buffer.BS_buffer\[68\] _3008_
+ _1179_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__a221oi_1
X_6134_ clknet_1_0__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__buf_1
X_3346_ BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__inv_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5016_ _1790_ _1792_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__nand3b_1
X_3277_ BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__inv_2
X_5918_ _2503_ _2516_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5849_ _2461_ _2471_ _2608_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__a21oi_2
X_6138__65 clknet_1_0__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__inv_2
XFILLER_0_86_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3200_ _2695_ _2711_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__nand2_2
X_4180_ BitStream_buffer.BS_buffer\[53\] _2986_ _2988_ BitStream_buffer.BS_buffer\[54\]
+ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__a22o_1
X_3131_ BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6080__12 clknet_1_0__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__inv_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ BitStream_buffer.BS_buffer\[57\] _2981_ _2983_ BitStream_buffer.BS_buffer\[58\]
+ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5703_ _2319_ _2327_ vssd1 vssd1 vccd1 vccd1 _2328_ sky130_fd_sc_hd__nor2_2
X_3895_ BitStream_buffer.BS_buffer\[73\] _2679_ _2682_ BitStream_buffer.BS_buffer\[74\]
+ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5634_ _2274_ _2261_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__and2_1
X_5981__82 clknet_1_0__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__inv_2
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ net1 BitStream_buffer.BS_buffer\[95\] _2192_ vssd1 vssd1 vccd1 vccd1 _2226_
+ sky130_fd_sc_hd__mux2_1
X_4516_ BitStream_buffer.BS_buffer\[28\] _0351_ _0380_ _0354_ _1299_ vssd1 vssd1 vccd1
+ vccd1 _1300_ sky130_fd_sc_hd__a221oi_1
X_5496_ _2178_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
X_4447_ _2765_ _2736_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__nand2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ _2956_ _2916_ _0847_ _2920_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__o22ai_1
X_3329_ _2862_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__buf_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3680_ _2859_ BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6117__46 clknet_1_1__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__inv_2
X_5350_ _0404_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__buf_2
X_5281_ net4 BitStream_buffer.BS_buffer\[35\] _2024_ vssd1 vssd1 vccd1 vccd1 _2031_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4301_ _1083_ _1084_ _1085_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__or4_1
X_4232_ _2746_ _2725_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4163_ _0473_ _2900_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__or2_1
X_4094_ BitStream_buffer.BS_buffer\[28\] _0337_ _0380_ _0341_ _0881_ vssd1 vssd1 vccd1
+ vccd1 _0882_ sky130_fd_sc_hd__a221oi_1
X_3114_ _2647_ _2642_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__nand2_4
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4996_ _0514_ _2848_ _1772_ _1773_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__o2111a_1
X_3947_ _2894_ _2890_ _0733_ _0734_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3878_ _0625_ _0637_ _0667_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5617_ _2262_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
X_5548_ _2214_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5479_ _2166_ _2148_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__and2_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _2742_ _2669_ _0686_ _2674_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3801_ _2775_ _2813_ _0588_ _0589_ _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__o2111a_1
X_4781_ _0468_ _2828_ _1559_ _1560_ _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__o2111a_1
X_3732_ BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3663_ _0453_ _2808_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5402_ _0405_ BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__nand2_1
X_5333_ _2067_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
X_3594_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5264_ net32 _2017_ _2018_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5195_ _1965_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_1
X_4215_ BitStream_buffer.BS_buffer\[80\] _2617_ BitStream_buffer.BS_buffer\[81\] _2624_
+ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__a221oi_1
X_4146_ _0444_ _2824_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__or2_1
X_4077_ BitStream_buffer.BS_buffer\[60\] _2992_ BitStream_buffer.BS_buffer\[61\] _2995_
+ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4979_ _0473_ _2779_ _1755_ _1756_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4000_ _2599_ _0786_ _0788_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__o21a_1
X_5951_ _2543_ _2542_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4902_ _0619_ _2908_ _0492_ _2911_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ _2404_ _2394_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__nand2_1
X_4833_ BitStream_buffer.BS_buffer\[27\] _0364_ BitStream_buffer.BS_buffer\[28\] _0368_
+ _1613_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__a221oi_1
X_4764_ _0453_ _2758_ _1542_ _1543_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3715_ _0505_ _2998_ _2996_ _3001_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__o22ai_1
X_4695_ BitStream_buffer.BS_buffer\[42\] _2928_ _2930_ BitStream_buffer.BS_buffer\[43\]
+ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__a22o_1
X_3646_ BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3577_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6296_ net98 _0311_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_5316_ _0404_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__buf_2
X_5247_ _2004_ _2005_ net30 _2001_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__a211o_1
X_5178_ net6 BitStream_buffer.BS_buffer\[1\] _1950_ vssd1 vssd1 vccd1 vccd1 _1954_
+ sky130_fd_sc_hd__mux2_1
X_4129_ _0437_ _2753_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3500_ _3033_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__buf_2
X_4480_ _1255_ _1257_ _1259_ _1263_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3431_ _2964_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__clkbuf_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ net112 _0165_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[126\] sky130_fd_sc_hd__dfxtp_2
X_3362_ _2895_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__clkbuf_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _0640_ _2848_ _1876_ _1877_ _1878_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__o2111a_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3293_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__inv_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ BitStream_buffer.BS_buffer\[25\] _3047_ _3049_ BitStream_buffer.BS_buffer\[26\]
+ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5934_ _2539_ _2549_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__nand2_1
X_5865_ _2485_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.exp_golomb_len\[1\] sky130_fd_sc_hd__inv_2
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4816_ _1592_ _1594_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5796_ _2307_ _2376_ _2378_ _2418_ _2420_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__a32o_1
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4747_ _1526_ _1527_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__nor2_1
X_4678_ _0638_ _2851_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__or2_1
X_3629_ _0419_ _2697_ _2694_ _2702_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__o22ai_1
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding_output[7] sky130_fd_sc_hd__buf_12
X_6279_ net81 _0294_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[12\] sky130_fd_sc_hd__dfxtp_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _3056_ _3062_ _0648_ _0323_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5650_ _2284_ _2285_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_0__f__2585_ clknet_0__2585_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2585_
+ sky130_fd_sc_hd__clkbuf_16
X_4601_ _1380_ _1381_ _1382_ _1383_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__or4_1
X_6023__121 clknet_1_1__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XFILLER_0_4_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _2237_ _2216_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4532_ _0407_ _2656_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4463_ _2831_ BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3414_ _2922_ _2634_ vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6202_ net164 _0217_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[74\] sky130_fd_sc_hd__dfxtp_2
X_4394_ _2664_ _3011_ BitStream_buffer.BS_buffer\[70\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _1179_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3345_ _2878_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__buf_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3276_ _2795_ _2797_ _2801_ _2805_ _2809_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__o2111a_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ BitStream_buffer.BS_buffer\[53\] _2948_ BitStream_buffer.BS_buffer\[54\] _2951_
+ _1793_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5917_ _2531_ _2533_ _2417_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _2464_ _2470_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__nor2_1
X_5779_ BitStream_buffer.BitStream_buffer_output\[8\] BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3130_ BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ _0499_ _2974_ _2963_ _2977_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5702_ _2317_ _2323_ _2326_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__a21o_1
X_3894_ _2631_ _2670_ _0556_ _2675_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5633_ net4 BitStream_buffer.BS_buffer\[115\] _2267_ vssd1 vssd1 vccd1 vccd1 _2274_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5564_ _2225_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
X_4515_ _0384_ _0357_ _0388_ _0360_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5495_ _2177_ _2171_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__and2_1
X_4446_ _2761_ BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__nand2_1
X_4377_ _0495_ _2909_ _2953_ _2912_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _2854_ _2677_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__nor2_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _2791_ _2792_ vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5280_ _2030_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
X_4300_ BitStream_buffer.BS_buffer\[15\] _0327_ _0329_ _0521_ vssd1 vssd1 vccd1 vccd1
+ _1086_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ _2820_ _2729_ BitStream_buffer.BS_buffer\[101\] _2732_ _1016_ vssd1 vssd1
+ vccd1 vccd1 _1017_ sky130_fd_sc_hd__a221oi_1
X_4162_ _0727_ _2896_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__or2_1
X_4093_ _0384_ _0344_ _0388_ _0347_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__o22ai_1
X_3113_ _2613_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4995_ _2858_ _3037_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__nand2_1
X_3946_ _2870_ _2900_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3877_ _0653_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5616_ _2260_ _2261_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__and2_1
X_5547_ _2213_ _2195_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__and2_1
X_5478_ net3 BitStream_buffer.BS_buffer\[68\] _2157_ vssd1 vssd1 vccd1 vccd1 _2166_
+ sky130_fd_sc_hd__mux2_1
X_4429_ _2631_ _2646_ _1210_ _1211_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__o2111a_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4780_ _0727_ _2840_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__or2_1
X_3800_ _2811_ _2824_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__or2_1
X_3731_ BitStream_buffer.BS_buffer\[13\] _3048_ _3050_ _0521_ vssd1 vssd1 vccd1 vccd1
+ _0522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3662_ _2804_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5401_ _2113_ _2098_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc\[2\] sky130_fd_sc_hd__xnor2_4
X_3593_ _2690_ _0338_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__nand2_2
X_5332_ _2066_ _2055_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6059__153 clknet_1_1__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
X_5263_ _2017_ net32 _0673_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5194_ _1964_ _1952_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__and2_1
X_4214_ _0560_ _2630_ _0419_ _2637_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4145_ _2819_ BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ _0508_ _2998_ _3009_ _3001_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4978_ _2790_ BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3929_ _2831_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5950_ _2512_ _2532_ _2557_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4901_ _1635_ _1650_ _1667_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5881_ BitStream_buffer.BitStream_buffer_output\[9\] _2466_ vssd1 vssd1 vccd1 vccd1
+ _2499_ sky130_fd_sc_hd__nor2_1
X_4832_ _0388_ _0371_ _0654_ _0374_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__o22ai_1
X_4763_ _0694_ _2770_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__or2_1
X_4694_ BitStream_buffer.BS_buffer\[48\] _2923_ _2925_ BitStream_buffer.BS_buffer\[49\]
+ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__a22o_1
X_3714_ BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3645_ _0431_ _2744_ _0432_ _0433_ _0435_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3576_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6295_ net97 _0310_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5315_ net8 BitStream_buffer.BS_buffer\[46\] _2023_ vssd1 vssd1 vccd1 vccd1 _2054_
+ sky130_fd_sc_hd__mux2_1
X_5246_ _1989_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5177_ _1953_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__clkbuf_1
X_4128_ _2749_ _2768_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__nand2_1
X_4059_ BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3430_ _2708_ BitStream_buffer.pc\[4\] BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1
+ vccd1 _2964_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3361_ _2659_ _2846_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__nand2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5100_ _2858_ _0516_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__nand2_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _1806_ _1807_ _1808_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__or4_1
X_6087__19 clknet_1_1__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__inv_2
X_3292_ _2811_ _2813_ _2817_ _2821_ _2825_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__o2111a_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5933_ _2548_ _2415_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__nand2_1
X_5988__89 clknet_1_1__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
X_5864_ _2608_ _2310_ _2353_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4815_ BitStream_buffer.BS_buffer\[71\] _3004_ BitStream_buffer.BS_buffer\[72\] _3007_
+ _1595_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5795_ _2419_ _2374_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4746_ BitStream_buffer.BS_buffer\[81\] _2678_ _2681_ BitStream_buffer.BS_buffer\[82\]
+ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4677_ _1446_ _1450_ _1454_ _1458_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3628_ BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
X_6000__100 clknet_1_1__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 half_fill_counter[0] sky130_fd_sc_hd__buf_12
X_3559_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__buf_2
X_6278_ net80 _0293_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[13\] sky130_fd_sc_hd__dfxtp_1
X_5229_ net28 _1988_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2584_ clknet_0__2584_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2584_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4600_ BitStream_buffer.BS_buffer\[57\] _2986_ _2988_ BitStream_buffer.BS_buffer\[58\]
+ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__a22o_1
X_5580_ net4 BitStream_buffer.BS_buffer\[99\] _2230_ vssd1 vssd1 vccd1 vccd1 _2237_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ _2650_ BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__nand2_1
X_4462_ _2827_ _2813_ _1243_ _1244_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3413_ BitStream_buffer.BS_buffer\[44\] _2935_ BitStream_buffer.BS_buffer\[45\] _2938_
+ _2946_ vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__a221oi_2
X_6201_ net163 _0216_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[75\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4393_ BitStream_buffer.BS_buffer\[63\] _2992_ BitStream_buffer.BS_buffer\[64\] _2995_
+ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a221oi_1
X_3344_ _2877_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__clkbuf_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _2806_ _2808_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__or2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _0750_ _2954_ _0626_ _2958_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__o22ai_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5916_ _2518_ _2519_ _2532_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5847_ _2348_ _2468_ _2442_ _2469_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__a22o_1
X_5778_ _2356_ _2353_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__nand2_1
X_4729_ _0847_ _0385_ _0739_ _0389_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6007__106 clknet_1_0__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6053__148 clknet_1_1__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_0_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5701_ _2324_ _2325_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__nand2_2
X_3962_ _0750_ _2967_ _0626_ _2970_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3893_ _2658_ _2646_ _0679_ _0680_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__o2111a_1
X_5632_ _2273_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5563_ _2224_ _2216_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__and2_1
X_4514_ BitStream_buffer.BS_buffer\[32\] _0337_ BitStream_buffer.BS_buffer\[33\] _0341_
+ _1297_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__a221oi_1
X_5494_ net13 BitStream_buffer.BS_buffer\[73\] _2157_ vssd1 vssd1 vccd1 vccd1 _2177_
+ sky130_fd_sc_hd__mux2_1
X_4445_ _2707_ _2744_ _1226_ _1227_ _1228_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__o2111a_1
X_6143__70 clknet_1_1__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__inv_2
X_4376_ _1115_ _1130_ _1147_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__and4_1
X_3327_ _2845_ _2849_ _2853_ _2857_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__o2111a_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__clkbuf_4
X_6046_ clknet_1_1__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__buf_1
X_3189_ _2710_ _2634_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4230_ _2795_ _2735_ _0453_ _2739_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__o22ai_1
X_4161_ _2892_ BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ _0874_ _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__nor2_1
X_3112_ _2645_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4994_ _2855_ BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__nand2_1
X_3945_ _0473_ _2896_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3876_ _0656_ _0659_ _0662_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__and4_1
X_5615_ net19 vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5546_ net13 _2706_ _2193_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__mux2_1
X_5477_ _2165_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
X_4428_ _0549_ _2661_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__or2_1
X_6036__132 clknet_1_0__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
X_4359_ _2835_ BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__nand2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6122__51 clknet_1_0__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__inv_2
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3730_ BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3661_ _2803_ BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3592_ BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
X_5400_ _2099_ _2100_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_42_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5331_ net5 BitStream_buffer.BS_buffer\[18\] _2061_ vssd1 vssd1 vccd1 vccd1 _2066_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5262_ _1986_ _1938_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4213_ _2599_ _0997_ _0999_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__o21a_1
X_5193_ net16 _0516_ _1950_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__mux2_1
X_4144_ _2815_ _2781_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4075_ _0859_ _0860_ _0861_ _0862_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4977_ _2786_ BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3928_ _0444_ _2813_ _0714_ _0715_ _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3859_ _0648_ _3062_ _0525_ _0323_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__o22ai_1
X_5529_ _2201_ _2195_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5880_ _1102_ _2467_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4900_ _1671_ _1673_ _1675_ _1679_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__and4_1
X_4831_ BitStream_buffer.BS_buffer\[32\] _0353_ BitStream_buffer.BS_buffer\[31\] _0351_
+ _1611_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4762_ _2764_ BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4693_ _0622_ _2915_ _0495_ _2919_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__o22ai_1
X_3713_ _0500_ _0501_ _0502_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__or4_1
X_3644_ _0434_ _2753_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3575_ _2654_ _0334_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6294_ net96 _0309_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5314_ _2053_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__clkbuf_1
X_5245_ _1988_ net28 vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__nand2_1
X_5176_ _1951_ _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__and2_1
X_4127_ _2746_ _2756_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4058_ _0800_ _0815_ _0832_ _0845_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3360_ BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__inv_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ BitStream_buffer.BS_buffer\[15\] _3040_ _3042_ _0363_ vssd1 vssd1 vccd1 vccd1
+ _1809_ sky130_fd_sc_hd__a22o_1
X_3291_ _2822_ _2824_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__or2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5932_ _2540_ _2547_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5863_ _2484_ vssd1 vssd1 vccd1 vccd1 exp_golomb_decoding.te_range\[2\] sky130_fd_sc_hd__inv_2
X_5794_ _2414_ _2607_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _2625_ _3010_ BitStream_buffer.BS_buffer\[74\] _3013_ vssd1 vssd1 vccd1 vccd1
+ _1595_ sky130_fd_sc_hd__a2bb2o_1
X_4745_ _0686_ _2669_ _0560_ _2674_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4676_ _2850_ _2828_ _1455_ _1456_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3627_ _0416_ _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__nor2_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 half_fill_counter[1] sky130_fd_sc_hd__buf_12
X_3558_ _0335_ _2672_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__nor2_2
X_6277_ net79 _0292_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[14\] sky130_fd_sc_hd__dfxtp_1
X_3489_ _3018_ _3022_ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__nor2_1
X_5228_ net29 vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__inv_2
X_5159_ net34 vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6092__23 clknet_1_1__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__inv_2
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2583_ clknet_0__2583_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2583_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5993__93 clknet_1_0__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
XFILLER_0_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4530_ BitStream_buffer.BS_buffer\[83\] _2617_ _2766_ _2624_ _1312_ vssd1 vssd1 vccd1
+ vccd1 _1313_ sky130_fd_sc_hd__a221oi_1
X_4461_ _2839_ _2824_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6200_ net162 _0215_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[76\] sky130_fd_sc_hd__dfxtp_2
X_3412_ _2939_ _2941_ _2942_ _2945_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4392_ _0411_ _2998_ _2652_ _3001_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3343_ _2690_ _2847_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__and2_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _2807_ vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__clkbuf_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ BitStream_buffer.BS_buffer\[57\] _2934_ BitStream_buffer.BS_buffer\[58\] _2937_
+ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__a221oi_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030__127 clknet_1_0__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
X_5915_ _2530_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__inv_2
X_5846_ BitStream_buffer.BitStream_buffer_output\[10\] _2397_ _2404_ vssd1 vssd1 vccd1
+ vccd1 _2469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5777_ BitStream_buffer.BitStream_buffer_output\[12\] BitStream_buffer.BitStream_buffer_output\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__xor2_1
X_4728_ BitStream_buffer.BS_buffer\[26\] _0364_ BitStream_buffer.BS_buffer\[27\] _0368_
+ _1509_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4659_ _2806_ _2758_ _1438_ _1439_ _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6129__57 clknet_1_0__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__inv_2
XFILLER_0_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5700_ BitStream_buffer.BitStream_buffer_output\[13\] BitStream_buffer.BitStream_buffer_output\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3892_ _0415_ _2661_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__or2_1
X_5631_ _2272_ _2261_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__and2_1
X_5562_ net8 BitStream_buffer.BS_buffer\[94\] _2192_ vssd1 vssd1 vccd1 vccd1 _2224_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4513_ _2914_ _0344_ _2917_ _0347_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__o22ai_1
X_5493_ _2176_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
X_4444_ _2715_ _2753_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__or2_1
X_4375_ _1151_ _1153_ _1155_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__and4_1
X_3326_ _2859_ BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__nand2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _2790_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__buf_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ _2720_ _2721_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5829_ _2451_ _2448_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__nand2_1
X_5972__74 clknet_1_1__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__inv_2
XFILLER_0_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4160_ _3044_ _2876_ _0518_ _2879_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__a221oi_1
X_3111_ _2644_ _2621_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__nand2_2
X_4091_ _0875_ _0876_ _0877_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4993_ _3027_ _2851_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__or2_1
X_3944_ _2892_ BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3875_ _0387_ _0379_ BitStream_buffer.BS_buffer\[31\] _0383_ _0664_ vssd1 vssd1 vccd1
+ vccd1 _0665_ sky130_fd_sc_hd__a221oi_1
X_5614_ net8 _2836_ _2229_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5545_ _2212_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6108__38 clknet_1_0__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__inv_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ _2164_ _2148_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__and2_1
X_4427_ _2625_ _2656_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__or2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _2831_ BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _2827_ _2829_ _2833_ _2837_ _2842_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__o2111a_1
X_4289_ _2671_ _3011_ BitStream_buffer.BS_buffer\[69\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _1075_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3660_ _2799_ BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3591_ _0382_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5330_ _2065_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5261_ _2015_ _2016_ _0675_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__a21oi_1
X_4212_ _0998_ _0672_ _0675_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__a21oi_1
X_5192_ _1963_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ _0456_ _2797_ _0927_ _0928_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__o2111a_1
X_4074_ BitStream_buffer.BS_buffer\[52\] _2986_ _2988_ BitStream_buffer.BS_buffer\[53\]
+ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4976_ _0727_ _2783_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__or2_1
X_3927_ _0456_ _2824_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3858_ BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3789_ _0567_ _0570_ _0574_ _0578_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__and4_1
X_5528_ net4 BitStream_buffer.BS_buffer\[83\] _2193_ vssd1 vssd1 vccd1 vccd1 _2201_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5459_ _2152_ _2148_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4830_ _2917_ _0356_ _0663_ _0359_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__o22ai_1
X_4761_ _2760_ BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4692_ _2939_ _2908_ _2942_ _2911_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__o22ai_1
X_3712_ BitStream_buffer.BS_buffer\[49\] _2986_ _2988_ BitStream_buffer.BS_buffer\[50\]
+ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3643_ BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3574_ BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__buf_2
X_5313_ _2052_ _2034_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__and2_1
X_6293_ net95 _0308_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_5244_ _2002_ _2003_ _0675_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__a21oi_1
X_5175_ _0404_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4126_ BitStream_buffer.BS_buffer\[99\] _2729_ _2820_ _2732_ _0912_ vssd1 vssd1 vccd1
+ vccd1 _0913_ sky130_fd_sc_hd__a221oi_1
X_4057_ _0836_ _0838_ _0840_ _0844_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _2714_ _2688_ _2736_ _2692_ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _2823_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__clkbuf_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5931_ _2545_ _2546_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__nand2_1
X_5862_ _2482_ _2307_ _2483_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5793_ _2375_ _2379_ _2416_ _2417_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__a22o_1
X_4813_ BitStream_buffer.BS_buffer\[67\] _2991_ BitStream_buffer.BS_buffer\[68\] _2994_
+ _1593_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4744_ _0549_ _2645_ _1522_ _1523_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4675_ _0601_ _2840_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__or2_1
X_3626_ BitStream_buffer.BS_buffer\[71\] _2679_ _2682_ BitStream_buffer.BS_buffer\[72\]
+ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__a22o_1
X_3557_ BitStream_buffer.BS_buffer\[24\] _0337_ BitStream_buffer.BS_buffer\[25\] _0341_
+ _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__a221oi_1
X_6276_ net78 _0291_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[15\] sky130_fd_sc_hd__dfxtp_2
X_5227_ _0403_ _1987_ _0405_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__o21ai_1
X_3488_ _3021_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__buf_4
X_5158_ _0672_ _1933_ _1935_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o21a_1
X_5089_ _2814_ BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__nand2_1
X_4109_ _0419_ _2630_ _2694_ _2637_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6077__10 clknet_1_0__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__inv_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5978__80 clknet_1_0__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__inv_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2582_ clknet_0__2582_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2582_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4460_ _2819_ _2832_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__nand2_1
X_3411_ _2944_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__buf_2
X_4391_ _1172_ _1173_ _1174_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or4_1
X_3342_ _2875_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__buf_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _2654_ _2778_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__nand2_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _0505_ _2940_ _2996_ _2944_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__o22ai_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5914_ _2520_ _2530_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__nand2_1
X_5845_ _2465_ _2467_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5776_ _2398_ _2400_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4727_ _0654_ _0371_ _0531_ _0374_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__o22ai_1
X_4658_ _0568_ _2770_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__or2_1
X_3609_ _0399_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__nand2_1
X_4589_ BitStream_buffer.BS_buffer\[47\] _2924_ _2926_ BitStream_buffer.BS_buffer\[48\]
+ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__a22o_1
X_6259_ net61 _0274_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[40\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ _0744_ _0746_ _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_57_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3891_ _2671_ _2656_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ net5 BitStream_buffer.BS_buffer\[114\] _2267_ vssd1 vssd1 vccd1 vccd1 _2272_
+ sky130_fd_sc_hd__mux2_1
X_5561_ _2223_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5492_ _2175_ _2171_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__and2_1
X_4512_ _1290_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4443_ _2749_ _2725_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4374_ _0601_ _2890_ _1156_ _1157_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__o2111a_1
X_3325_ _2858_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__buf_4
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _2777_ _2634_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__nor2_2
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5828_ _2449_ _2375_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5759_ _2370_ _2383_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ _2643_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4090_ _3051_ _0327_ _0329_ _0770_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4992_ _1758_ _1762_ _1766_ _1770_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3943_ BitStream_buffer.BS_buffer\[1\] _2876_ _3039_ _2879_ _0731_ vssd1 vssd1 vccd1
+ vccd1 _0732_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3874_ _0663_ _0386_ _0540_ _0390_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__o22ai_1
X_5613_ _2259_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
X_5544_ _2211_ _2195_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__and2_1
X_5475_ net4 BitStream_buffer.BS_buffer\[67\] _2157_ vssd1 vssd1 vccd1 vccd1 _2164_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4426_ _2650_ BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nand2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _0464_ _2813_ _1139_ _1140_ _1141_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__o2111a_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _2839_ _2841_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__or2_1
X_4288_ BitStream_buffer.BS_buffer\[62\] _2992_ BitStream_buffer.BS_buffer\[63\] _2995_
+ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__a221oi_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _2757_ _2759_ _2763_ _2767_ _2772_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_64_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5260_ net34 net33 vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__nand2_1
X_4211_ BitStream_buffer.BitStream_buffer_output\[10\] vssd1 vssd1 vccd1 vccd1 _0998_
+ sky130_fd_sc_hd__inv_2
X_6113__42 clknet_1_1__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__inv_2
X_5191_ _1962_ _1952_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__and2_1
X_4142_ _0459_ _2808_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__or2_1
X_4073_ BitStream_buffer.BS_buffer\[58\] _2981_ _2983_ BitStream_buffer.BS_buffer\[59\]
+ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ _1743_ _1745_ _1749_ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__and4_1
X_3926_ _2819_ BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3857_ _0646_ _3055_ _0523_ _3058_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3788_ _2707_ _2759_ _0575_ _0576_ _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__o2111a_1
X_5527_ _2200_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5458_ net8 BitStream_buffer.BS_buffer\[62\] _2120_ vssd1 vssd1 vccd1 vccd1 _2152_
+ sky130_fd_sc_hd__mux2_1
X_5389_ _2107_ _2105_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc\[5\] sky130_fd_sc_hd__nor2_2
X_4409_ BitStream_buffer.BS_buffer\[32\] _0340_ BitStream_buffer.BS_buffer\[31\] _0337_
+ _1193_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_5_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4760_ _2737_ _2743_ _1538_ _1539_ _1540_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__o2111a_1
X_4691_ _1427_ _1442_ _1459_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__and4_1
X_3711_ BitStream_buffer.BS_buffer\[55\] _2981_ _2983_ BitStream_buffer.BS_buffer\[56\]
+ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3642_ _2749_ BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3573_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__buf_2
X_5312_ net9 BitStream_buffer.BS_buffer\[45\] _2023_ vssd1 vssd1 vccd1 vccd1 _2052_
+ sky130_fd_sc_hd__mux2_1
X_6292_ net94 _0307_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5243_ _2001_ net30 vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__nand2_1
X_5174_ net7 _0400_ _1950_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__mux2_1
X_4125_ _0453_ _2735_ _2806_ _2739_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4056_ _2870_ _2890_ _0841_ _0842_ _0843_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4958_ _0423_ _2696_ _2707_ _2701_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__o22ai_1
X_4889_ _2855_ _0516_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__nand2_1
X_3909_ _2749_ BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6049__144 clknet_1_0__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
XFILLER_0_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5930_ _2489_ _2541_ _2543_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5861_ _2478_ _2480_ _2479_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__nand3_1
X_5792_ net17 _2605_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__nor2_2
X_4812_ _0415_ _2997_ _2664_ _3000_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4743_ _0419_ _2660_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4674_ _2834_ BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__nand2_1
X_3625_ _0415_ _2670_ _2664_ _2675_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__o22ai_1
X_3556_ _0342_ _0344_ _0345_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6275_ net77 _0290_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_valid_n
+ sky130_fd_sc_hd__dfxtp_1
X_5226_ _1985_ net32 _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__and3_1
X_3487_ _2654_ _3020_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__nand2_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5157_ _1934_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__a21oi_1
X_4108_ _2599_ _0893_ _0895_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__o21a_1
X_5088_ _2898_ _2796_ _1863_ _1864_ _1865_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__o2111a_1
X_4039_ _2782_ _2813_ _0824_ _0825_ _0826_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__2581_ clknet_0__2581_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2581_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3410_ _2943_ _2907_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__nand2_2
X_4390_ BitStream_buffer.BS_buffer\[55\] _2986_ _2988_ BitStream_buffer.BS_buffer\[56\]
+ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3341_ _2854_ _2687_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__nor2_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__inv_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _1786_ _1787_ _1788_ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__or4_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5913_ _2529_ _2415_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__nand2_1
X_5844_ _2466_ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5775_ _2363_ _2326_ _2399_ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__nand3_1
XFILLER_0_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4726_ _0387_ _0350_ BitStream_buffer.BS_buffer\[31\] _0353_ _1507_ vssd1 vssd1 vccd1
+ vccd1 _1508_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4657_ _2764_ BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3608_ BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4588_ _0495_ _2916_ _2953_ _2920_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__o22ai_1
X_3539_ _0325_ _0327_ _0329_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__a22o_1
X_6258_ net60 _0273_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[41\] sky130_fd_sc_hd__dfxtp_2
X_6189_ net151 _0204_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[87\] sky130_fd_sc_hd__dfxtp_1
X_5209_ net11 _0650_ _1949_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3890_ _2650_ BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__nand2_1
X_5560_ _2222_ _2216_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4511_ _1291_ _1292_ _1293_ _1294_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5491_ net14 BitStream_buffer.BS_buffer\[72\] _2157_ vssd1 vssd1 vccd1 vccd1 _2175_
+ sky130_fd_sc_hd__mux2_1
X_4442_ _2746_ _2721_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__nand2_1
X_4373_ _0727_ _2900_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__or2_1
X_6112_ clknet_1_0__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__buf_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _2854_ _2634_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__nor2_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _2787_ _2788_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__nand2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _2719_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5827_ _2419_ _2421_ _2450_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__o21ai_2
X_5758_ _2380_ _2382_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__nand2_1
X_4709_ _2631_ _3010_ BitStream_buffer.BS_buffer\[73\] _3013_ vssd1 vssd1 vccd1 vccd1
+ _1491_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5689_ BitStream_buffer.BitStream_buffer_output\[13\] _2313_ vssd1 vssd1 vccd1 vccd1
+ _2314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4991_ _2883_ _2828_ _1767_ _1768_ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _0730_ _2882_ _0604_ _2885_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3873_ BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5612_ _2258_ _2240_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__and2_1
X_5543_ net14 _2725_ _2193_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5474_ _2163_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
X_4425_ BitStream_buffer.BS_buffer\[82\] _2617_ BitStream_buffer.BS_buffer\[83\] _2624_
+ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4356_ _0445_ _2824_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__or2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _2840_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__clkbuf_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _2652_ _2998_ _2640_ _3001_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__o22ai_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _2769_ _2771_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__or2_1
X_3169_ _2694_ _2697_ _2698_ _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6043__139 clknet_1_1__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ _0953_ _0995_ _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__nand3_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5190_ net2 _3037_ _1950_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__mux2_1
X_4141_ _2803_ BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nand2_1
X_4072_ _0626_ _2974_ _0499_ _2977_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__o22ai_1
X_4974_ _0450_ _2758_ _1750_ _1751_ _1752_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__o2111a_1
X_3925_ _2815_ BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3856_ BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3787_ _2757_ _2771_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or2_1
X_5526_ _2199_ _2195_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__and2_1
X_5457_ _2151_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
X_4408_ _2917_ _0344_ _0663_ _0347_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5388_ _2104_ BitStream_buffer.pc_previous\[4\] BitStream_buffer.pc_previous\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4339_ _0423_ _2753_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6026__123 clknet_1_0__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
X_3710_ _2968_ _2974_ _2972_ _2977_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__o22ai_1
X_4690_ _1463_ _1465_ _1467_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3641_ _2746_ BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3572_ _0335_ _2643_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5311_ _2051_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__clkbuf_1
X_6291_ net93 _0306_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5242_ net30 net28 _1940_ _1989_ _2001_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__a2111o_1
X_5173_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__clkbuf_4
X_4124_ _0428_ _2713_ _0908_ _0909_ _0910_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__o2111a_1
Xinput1 BitStream_buffer_input[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
X_4055_ _2867_ _2900_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4957_ _1734_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__nor2_1
X_4888_ _0869_ _2851_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3908_ _2746_ _2768_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__nand2_1
X_3839_ BitStream_buffer.BS_buffer\[56\] _2981_ _2983_ BitStream_buffer.BS_buffer\[57\]
+ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5509_ net8 BitStream_buffer.BS_buffer\[78\] _2156_ vssd1 vssd1 vccd1 vccd1 _2187_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5860_ net22 _2481_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4811_ _1588_ _1589_ _1590_ _1591_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5791_ _2414_ _2415_ _2373_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4742_ _2698_ _2655_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4673_ _2830_ BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3624_ BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3555_ _0346_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6274_ net76 _0289_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dfxtp_2
X_3486_ _3019_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__clkbuf_4
X_5225_ net31 vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__inv_2
X_5156_ BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1 vccd1 _1934_
+ sky130_fd_sc_hd__inv_2
X_4107_ _0894_ _0672_ _0675_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__a21oi_1
X_5087_ _2827_ _2807_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__or2_1
X_4038_ _2775_ _2824_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2580_ clknet_0__2580_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2580_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3340_ BitStream_buffer.BS_buffer\[118\] _2863_ BitStream_buffer.BS_buffer\[119\]
+ _2866_ _2873_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__a221oi_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ BitStream_buffer.BS_buffer\[45\] _2928_ _2930_ BitStream_buffer.BS_buffer\[46\]
+ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a22o_1
X_3271_ _2803_ _2804_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__nand2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083__15 clknet_1_0__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__inv_2
X_5912_ _2526_ _2528_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5843_ _2321_ _2405_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5774_ BitStream_buffer.BitStream_buffer_output\[14\] BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__xnor2_1
X_5984__85 clknet_1_0__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__inv_2
X_4725_ _0663_ _0356_ _0540_ _0359_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4656_ _2760_ _2800_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__nand2_1
X_4587_ _2942_ _2909_ _0622_ _2912_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__o22ai_1
X_3607_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__buf_2
X_3538_ BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6257_ net59 _0272_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[42\] sky130_fd_sc_hd__dfxtp_2
X_3469_ BitStream_buffer.BS_buffer\[56\] _2992_ BitStream_buffer.BS_buffer\[57\] _2995_
+ _3002_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__a221oi_1
X_6188_ net150 _0203_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[88\] sky130_fd_sc_hd__dfxtp_1
X_5208_ _1974_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__clkbuf_1
X_5139_ _0657_ _3061_ _0534_ _0322_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5490_ _2174_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4510_ _0366_ _0327_ _0329_ _0363_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4441_ _2816_ _2729_ BitStream_buffer.BS_buffer\[103\] _2732_ _1224_ vssd1 vssd1
+ vccd1 vccd1 _1225_ sky130_fd_sc_hd__a221oi_1
X_4372_ _0468_ _2896_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__or2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _2856_ BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__nand2_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__clkbuf_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _2710_ _2615_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5826_ _2448_ _2417_ _2449_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5757_ _2381_ BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1 vccd1
+ _2382_ sky130_fd_sc_hd__nand2_1
X_4708_ BitStream_buffer.BS_buffer\[66\] _2991_ BitStream_buffer.BS_buffer\[67\] _2994_
+ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5688_ _0787_ _0894_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__nand2_1
X_4639_ _0407_ _2645_ _1418_ _1419_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6020__118 clknet_1_1__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4990_ _0468_ _2840_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3941_ _0400_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__inv_2
X_3872_ BitStream_buffer.BS_buffer\[18\] _0365_ BitStream_buffer.BS_buffer\[19\] _0369_
+ _0661_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5611_ net9 _2838_ _2229_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__mux2_1
X_5542_ _2210_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5473_ _2162_ _2148_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4424_ _2742_ _2630_ _0686_ _2637_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4355_ _2819_ _2781_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__nand2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _2695_ _2778_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__nand2_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _1068_ _1069_ _1070_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__or4_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _2770_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__clkbuf_2
X_3168_ _2701_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__buf_2
X_3099_ BitStream_buffer.pc\[2\] _2604_ _2632_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5809_ _0894_ _2394_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4140_ _2799_ BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__nand2_1
X_4071_ _0858_ _2967_ _0750_ _2970_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__o22ai_1
X_4973_ _0453_ _2770_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__or2_1
X_3924_ _0459_ _2797_ _0710_ _0711_ _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3855_ _0521_ _3048_ _3050_ BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1
+ _0645_ sky130_fd_sc_hd__a22o_1
X_3786_ _2765_ _2762_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__nand2_1
X_6003__102 clknet_1_0__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
XFILLER_0_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5525_ net5 BitStream_buffer.BS_buffer\[82\] _2193_ vssd1 vssd1 vccd1 vccd1 _2199_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ _2150_ _2148_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__and2_1
X_4407_ _1186_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__nor2_1
X_5387_ _2106_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__inv_2
X_4338_ _2749_ _2756_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_1
X_4269_ _0473_ _2890_ _1052_ _1053_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2597_ clknet_0__2597_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2597_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3640_ BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3571_ BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__buf_2
X_6290_ net92 _0305_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[1\] sky130_fd_sc_hd__dfxtp_2
X_5310_ _2050_ _2034_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5241_ _2000_ _1987_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__nand2_2
X_5172_ _1944_ _1948_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__nand2_4
X_4123_ _2724_ BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__nand2_1
Xinput2 BitStream_buffer_input[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_4
X_4054_ _0601_ _2896_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ BitStream_buffer.BS_buffer\[83\] _2678_ _2681_ _2766_ vssd1 vssd1 vccd1 vccd1
+ _1735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4887_ _1654_ _1658_ _1662_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__and4_1
X_3907_ BitStream_buffer.BS_buffer\[97\] _2729_ _2804_ _2732_ _0695_ vssd1 vssd1 vccd1
+ vccd1 _0696_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_34_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3838_ _2963_ _2974_ _2968_ _2977_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5508_ _2186_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
X_3769_ _0557_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__nor2_1
X_6089__21 clknet_1_1__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__inv_2
X_5439_ net14 BitStream_buffer.BS_buffer\[56\] _2121_ vssd1 vssd1 vccd1 vccd1 _2139_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4810_ BitStream_buffer.BS_buffer\[59\] _2985_ _2987_ BitStream_buffer.BS_buffer\[60\]
+ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__a22o_1
X_5790_ _2607_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4741_ _2649_ BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4672_ _2898_ _2812_ _1451_ _1452_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3623_ _2652_ _2646_ _0410_ _0412_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_24_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3554_ _2957_ _0338_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6273_ net75 _0288_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dfxtp_2
X_3485_ _2708_ _2600_ _2601_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__and3_1
X_5224_ net33 _1936_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__nor2_1
X_5155_ _1889_ _1931_ _1932_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4106_ BitStream_buffer.BitStream_buffer_output\[11\] vssd1 vssd1 vccd1 vccd1 _0894_
+ sky130_fd_sc_hd__inv_4
X_5086_ _2802_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _2819_ _2792_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4939_ _2953_ _0385_ _2956_ _0389_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6055__150 clknet_1_1__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3270_ BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__clkbuf_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5911_ _0998_ _2467_ _2527_ _2349_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5842_ _1206_ _2322_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5773_ _2393_ _2397_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__nand2_1
X_4724_ BitStream_buffer.BS_buffer\[34\] _0336_ BitStream_buffer.BS_buffer\[35\] _0341_
+ _1505_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4655_ _2715_ _2743_ _1434_ _1435_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3606_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__clkbuf_2
X_4586_ _1323_ _1338_ _1355_ _1368_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__and4_1
X_3537_ _0328_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__buf_2
X_6256_ net58 _0271_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[43\] sky130_fd_sc_hd__dfxtp_2
X_3468_ _2996_ _2998_ _2999_ _3001_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__o22ai_1
X_6187_ net149 _0202_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[89\] sky130_fd_sc_hd__dfxtp_1
X_5207_ _1972_ _1973_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__and2_1
X_3399_ _2913_ _2921_ _2927_ _2932_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__or4_1
X_5138_ _0654_ _3054_ _0531_ _3057_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__o22ai_1
X_5069_ _2811_ _2712_ _1844_ _1845_ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4440_ _2822_ _2735_ _0450_ _2739_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__o22ai_1
X_4371_ _2892_ BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__nand2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__buf_4
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _2786_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__buf_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _2715_ _2717_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5825_ _2446_ _2415_ _2414_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5756_ _2368_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__buf_6
XFILLER_0_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5687_ _2311_ _0403_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4707_ _2664_ _2997_ _2671_ _3000_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__o22ai_1
X_4638_ _2694_ _2660_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__or2_1
X_4569_ _2835_ BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nand2_1
X_6239_ net41 _0254_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[28\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6125__53 clknet_1_1__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__inv_2
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6140__67 clknet_1_1__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__inv_2
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3940_ BitStream_buffer.BS_buffer\[121\] _2863_ BitStream_buffer.BS_buffer\[122\]
+ _2866_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_58_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3871_ _0660_ _0372_ _0537_ _0375_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__o22ai_1
X_5610_ _2257_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
X_5541_ _2209_ _2195_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5472_ net5 BitStream_buffer.BS_buffer\[66\] _2157_ vssd1 vssd1 vccd1 vccd1 _2162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4423_ _2599_ _1205_ _1207_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__o21a_1
X_4354_ _2815_ _2838_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nand2_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3305_ _2838_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ BitStream_buffer.BS_buffer\[54\] _2986_ _2988_ BitStream_buffer.BS_buffer\[55\]
+ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__a22o_1
X_6024_ clknet_1_1__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__buf_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _2668_ _2711_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__nand2_1
X_3167_ _2700_ _2621_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3098_ _2612_ _2626_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5808_ BitStream_buffer.BitStream_buffer_output\[11\] _2395_ vssd1 vssd1 vccd1 vccd1
+ _2432_ sky130_fd_sc_hd__nor2_1
X_5739_ _2363_ _0671_ _2326_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4070_ BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__inv_2
X_4972_ _2764_ BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3923_ _0450_ _2808_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3854_ _0639_ _0641_ _0642_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3785_ _2761_ _2725_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__nand2_1
X_5524_ _2198_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5455_ net9 BitStream_buffer.BS_buffer\[61\] _2120_ vssd1 vssd1 vccd1 vccd1 _2150_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4406_ _1187_ _1188_ _1189_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__or4_1
X_5386_ _0405_ BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__nand2_1
X_6104__34 clknet_1_1__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__inv_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _2746_ _2706_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__nand2_1
X_4268_ _0601_ _2900_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__or2_1
X_3219_ _2752_ vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__clkbuf_2
X_4199_ _0380_ _0337_ _0387_ _0341_ _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2596_ clknet_0__2596_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2596_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ BitStream_buffer.BS_buffer\[20\] _0351_ BitStream_buffer.BS_buffer\[21\] _0354_
+ _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _1993_ _1998_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__nand3_1
X_5171_ _1945_ _1946_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__and3_1
X_4122_ _2720_ BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__nand2_1
X_4053_ _2892_ BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__nand2_1
Xinput3 BitStream_buffer_input[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_4
XFILLER_0_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4955_ _0431_ _2669_ _2742_ _2674_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__o22ai_1
X_3906_ _0694_ _2735_ _0568_ _2739_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__o22ai_1
X_4886_ _2845_ _2828_ _1663_ _1664_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3837_ _0626_ _2967_ _0499_ _2970_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3768_ BitStream_buffer.BS_buffer\[72\] _2679_ _2682_ BitStream_buffer.BS_buffer\[73\]
+ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__a22o_1
X_5507_ _2185_ _2171_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3699_ BitStream_buffer.BS_buffer\[33\] _2929_ _2931_ BitStream_buffer.BS_buffer\[34\]
+ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__a22o_1
X_5438_ _2138_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
X_5369_ _2091_ _2079_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4740_ _2768_ _2616_ _2762_ _2623_ _1520_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4671_ _2827_ _2823_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3622_ _2671_ _2661_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__or2_1
X_3553_ BitStream_buffer.BS_buffer\[26\] vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
X_6272_ net74 _0287_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dfxtp_2
X_3484_ BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__inv_2
X_5223_ _1984_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
X_5154_ _0398_ _0521_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__nand2_1
X_4105_ _0846_ _0891_ _0892_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__nand3_1
X_5085_ _2798_ _2836_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4036_ _2815_ _2788_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4938_ BitStream_buffer.BS_buffer\[28\] _0364_ _0380_ _0368_ _1717_ vssd1 vssd1 vccd1
+ vccd1 _1718_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_30 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4869_ _2795_ _2758_ _1646_ _1647_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5910_ _2397_ _2467_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5841_ _2393_ _2462_ _2463_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5772_ _2395_ _2396_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__nand2_1
X_4723_ _2905_ _0343_ _2910_ _0346_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4654_ _2733_ _2752_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__or2_1
X_4585_ _1359_ _1361_ _1363_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__and4_1
X_3605_ _0396_ _2708_ _2600_ _2601_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__and4_1
X_3536_ _3032_ _2634_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nor2_2
X_6039__135 clknet_1_0__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
X_6255_ net57 _0270_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[44\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5206_ _0404_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__buf_2
X_3467_ _3000_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__buf_2
X_6186_ net148 _0201_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[90\] sky130_fd_sc_hd__dfxtp_1
X_3398_ BitStream_buffer.BS_buffer\[32\] _2929_ _2931_ BitStream_buffer.BS_buffer\[33\]
+ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__a22o_1
X_5137_ BitStream_buffer.BS_buffer\[26\] _3047_ _3049_ BitStream_buffer.BS_buffer\[27\]
+ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__a22o_1
X_5068_ _2723_ _2816_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__nand2_1
X_4019_ _2746_ _2762_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4370_ _3037_ _2876_ _0516_ _2879_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__a221oi_1
X_3321_ _2854_ _2615_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _2777_ _2615_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__nor2_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _2716_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5824_ _2447_ _2419_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ _2366_ BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1 vccd1
+ _2380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5686_ BitStream_buffer.BitStream_buffer_output\[15\] BitStream_buffer.BitStream_buffer_output\[14\]
+ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__nor2_1
X_4706_ _1484_ _1485_ _1486_ _1487_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4637_ _0549_ _2655_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4568_ _2831_ BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__nand2_1
X_3519_ BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__inv_2
X_4499_ _0415_ _3011_ BitStream_buffer.BS_buffer\[71\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _1283_ sky130_fd_sc_hd__a2bb2o_1
X_6238_ net40 _0253_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[29\] sky130_fd_sc_hd__dfxtp_1
X_6169_ net131 _0184_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[107\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3870_ BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5540_ net15 _2756_ _2193_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__mux2_1
X_5471_ _2161_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4422_ _1206_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4353_ _0444_ _2797_ _1135_ _1136_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__o2111a_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__clkbuf_4
X_4284_ BitStream_buffer.BS_buffer\[60\] _2981_ _2983_ BitStream_buffer.BS_buffer\[61\]
+ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__a22o_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _2768_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__inv_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _2699_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__inv_2
X_3097_ BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3999_ _0787_ _0672_ _0675_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__a21oi_1
X_5807_ _2426_ _2430_ _2371_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__nand3_1
X_5738_ _2347_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _2298_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4971_ _2760_ BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__nand2_1
X_3922_ _2803_ BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__nand2_1
X_3853_ _0518_ _3041_ _3043_ _3037_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3784_ _2751_ _2744_ _0571_ _0572_ _0573_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_54_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5523_ _2197_ _2195_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5454_ _2149_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
X_5385_ BitStream_buffer.pc_previous\[6\] _2105_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc\[6\]
+ sky130_fd_sc_hd__xor2_4
X_4405_ _0363_ _0327_ _0329_ BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1
+ _1190_ sky130_fd_sc_hd__a22o_1
X_4336_ BitStream_buffer.BS_buffer\[101\] _2729_ _2816_ _2732_ _1120_ vssd1 vssd1
+ vccd1 vccd1 _1121_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_5_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4267_ _2850_ _2896_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__or2_1
X_4198_ _0540_ _0344_ _0384_ _0347_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__o22ai_1
X_3218_ _2659_ _2711_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__nand2_1
X_3149_ BitStream_buffer.BS_buffer\[70\] _2679_ _2682_ BitStream_buffer.BS_buffer\[71\]
+ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2595_ clknet_0__2595_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2595_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5170_ BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__inv_2
X_4121_ _0694_ _2717_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__or2_1
X_4052_ _3039_ _2876_ _3044_ _2879_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__a221oi_1
Xinput4 BitStream_buffer_input[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_4
X_4954_ _2694_ _2645_ _1730_ _1731_ _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_86_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3905_ _2800_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__inv_2
X_4885_ _2850_ _2840_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3767_ _0556_ _2670_ _0415_ _2675_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__o22ai_1
X_5506_ net9 BitStream_buffer.BS_buffer\[77\] _2156_ vssd1 vssd1 vccd1 vccd1 _2185_
+ sky130_fd_sc_hd__mux2_1
X_3698_ BitStream_buffer.BS_buffer\[39\] _2924_ _2926_ BitStream_buffer.BS_buffer\[40\]
+ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__a22o_1
X_5437_ _2137_ _2127_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5368_ net8 _0387_ _2060_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__mux2_1
X_5299_ _2043_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
X_4319_ _0686_ _2630_ _0560_ _2637_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_69_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095__26 clknet_1_0__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__inv_2
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5996__96 clknet_1_1__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
XFILLER_0_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4670_ _2818_ _2836_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__nand2_1
X_3621_ _0411_ _2656_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__or2_1
X_3552_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6271_ net73 _0286_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dfxtp_2
X_3483_ _2990_ _3003_ _3016_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__nand3b_1
X_5222_ _1983_ _1973_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5153_ _1899_ _1909_ _1930_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__nor3_1
X_4104_ _0399_ _0518_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nand2_1
X_5084_ _0601_ _2779_ _1859_ _1860_ _1861_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__o2111a_1
X_4035_ _2811_ _2797_ _0820_ _0821_ _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4937_ _0384_ _0371_ _0388_ _0374_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4868_ _2806_ _2770_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3819_ _2894_ _2900_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4799_ BitStream_buffer.BS_buffer\[49\] _2923_ _2925_ BitStream_buffer.BS_buffer\[50\]
+ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__a22o_1
Xclkbuf_0__2597_ _2597_ vssd1 vssd1 vccd1 vccd1 clknet_0__2597_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6016__114 clknet_1_0__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6062__156 clknet_1_0__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5840_ _2432_ BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1 vccd1 vccd1
+ _2463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5771_ BitStream_buffer.BitStream_buffer_output\[10\] BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4722_ _1498_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4653_ _2748_ _2721_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__nand2_1
X_4584_ _2850_ _2890_ _1364_ _1365_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__o2111a_1
X_3604_ _2612_ _2665_ _2604_ _2626_ _3032_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__a41o_1
XFILLER_0_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3535_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6254_ net56 _0269_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[45\] sky130_fd_sc_hd__dfxtp_2
X_3466_ _2957_ _2965_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__nand2_2
X_5205_ net12 _0527_ _1949_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__mux2_1
X_6185_ net147 _0200_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[91\] sky130_fd_sc_hd__dfxtp_1
X_3397_ _2930_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5136_ _1910_ _1911_ _1912_ _1913_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__or4_1
X_5067_ _2719_ _2792_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__nand2_1
X_4018_ _2804_ _2729_ BitStream_buffer.BS_buffer\[99\] _2732_ _0805_ vssd1 vssd1 vccd1
+ vccd1 _0806_ sky130_fd_sc_hd__a221oi_1
X_5969_ clknet_1_0__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__buf_1
X_5975__77 clknet_1_0__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__inv_2
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3320_ _2846_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__inv_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _2782_ _2784_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__or2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _2620_ _2711_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5823_ _2446_ _2415_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ net18 _2606_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5685_ _2308_ _2309_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__and2_2
X_4705_ BitStream_buffer.BS_buffer\[58\] _2985_ _2987_ BitStream_buffer.BS_buffer\[59\]
+ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4636_ _2649_ BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6306_ net37 _0321_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_4567_ _2888_ _2813_ _1347_ _1348_ _1349_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3518_ BitStream_buffer.BS_buffer\[12\] _3048_ _3050_ _3051_ vssd1 vssd1 vccd1 vccd1
+ _3052_ sky130_fd_sc_hd__a22o_1
X_4498_ BitStream_buffer.BS_buffer\[64\] _2992_ BitStream_buffer.BS_buffer\[65\] _2995_
+ _1281_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a221oi_1
X_6237_ net39 _0252_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[30\] sky130_fd_sc_hd__dfxtp_1
X_3449_ _2982_ vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__clkbuf_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ net130 _0183_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[108\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5119_ _0858_ _2954_ _0750_ _2958_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5470_ _2160_ _2148_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__and2_1
X_4421_ BitStream_buffer.BitStream_buffer_output\[8\] vssd1 vssd1 vccd1 vccd1 _1206_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ _0456_ _2808_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__or2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _2835_ _2836_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__nand2_1
X_4283_ _0858_ _2974_ _0750_ _2977_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__o22ai_1
X_3234_ BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__clkbuf_4
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _2641_ _2686_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__nand2_4
X_3096_ _2629_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6072__5 clknet_1_1__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__inv_2
X_3998_ BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1 vccd1 vccd1 _0787_
+ sky130_fd_sc_hd__inv_2
X_5806_ _2370_ _2429_ _2390_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__nand3_1
X_5737_ _2361_ _1102_ _2326_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5668_ _2297_ _2285_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4619_ BitStream_buffer.BS_buffer\[33\] _0337_ BitStream_buffer.BS_buffer\[34\] _0341_
+ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5599_ net13 BitStream_buffer.BS_buffer\[105\] _2230_ vssd1 vssd1 vccd1 vccd1 _2250_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _0428_ _2743_ _1746_ _1747_ _1748_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__o2111a_1
X_3921_ _2799_ BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3852_ _0516_ _3034_ _3036_ BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1
+ _0642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5522_ net6 BitStream_buffer.BS_buffer\[81\] _2193_ vssd1 vssd1 vccd1 vccd1 _2197_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3783_ _2769_ _2753_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5453_ _2147_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__and2_1
X_5384_ _2104_ BitStream_buffer.pc_previous\[4\] BitStream_buffer.pc_previous\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__and3_2
X_4404_ _0373_ _3062_ _0646_ _0323_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__o22ai_1
X_4335_ _0450_ _2735_ _2795_ _2739_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4266_ _2892_ BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4197_ _0978_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__nor2_1
X_3217_ BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__inv_2
X_6010__109 clknet_1_1__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
X_3148_ _2681_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__clkbuf_4
X_3079_ _2612_ BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2594_ clknet_0__2594_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2594_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4120_ _0897_ _0901_ _0904_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__and4_1
X_4051_ _3018_ _2882_ _0730_ _2885_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__o22ai_1
Xinput5 BitStream_buffer_input[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _0686_ _2660_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3904_ _2737_ _2713_ _0690_ _0691_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o2111a_1
X_4884_ _2834_ BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ _0618_ _0621_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__nand3b_1
X_3766_ BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5505_ _2184_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3697_ _2910_ _2916_ _2914_ _2920_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5436_ net15 BitStream_buffer.BS_buffer\[55\] _2121_ vssd1 vssd1 vccd1 vccd1 _2137_
+ sky130_fd_sc_hd__mux2_1
X_5367_ _2090_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4318_ _2599_ _1101_ _1103_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__o21a_1
X_5298_ _2042_ _2034_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__and2_1
X_4249_ _2815_ _2832_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3620_ BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3551_ net36 _0338_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__nand2_2
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ net72 _0285_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dfxtp_2
X_3482_ BitStream_buffer.BS_buffer\[60\] _3005_ BitStream_buffer.BS_buffer\[61\] _3008_
+ _3015_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__a221oi_1
X_5221_ net1 BitStream_buffer.BS_buffer\[15\] _1949_ vssd1 vssd1 vccd1 vccd1 _1983_
+ sky130_fd_sc_hd__mux2_1
X_5152_ _1920_ _1929_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__nand2_1
X_4103_ _0857_ _0868_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5083_ _2790_ BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4034_ _2822_ _2808_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4936_ BitStream_buffer.BS_buffer\[32\] _0350_ BitStream_buffer.BS_buffer\[33\] _0353_
+ _1715_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__a221oi_1
XANTENNA_10 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _1411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _2764_ _2800_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3818_ _2867_ _2896_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4798_ _2942_ _2915_ _0622_ _2919_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__o22ai_1
X_3749_ BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__inv_2
Xclkbuf_0__2596_ _2596_ vssd1 vssd1 vccd1 vccd1 clknet_0__2596_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5419_ _2125_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5770_ _2394_ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__inv_2
X_4721_ _1499_ _1500_ _1501_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4652_ _2745_ _2736_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__nand2_1
X_3603_ _2962_ _3017_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__nor3_1
X_4583_ _0468_ _2900_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3534_ _2628_ _3020_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__and2_2
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6253_ net55 _0268_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[46\] sky130_fd_sc_hd__dfxtp_2
X_3465_ BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__inv_2
X_5204_ _1971_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__clkbuf_1
X_6184_ net146 _0199_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[92\] sky130_fd_sc_hd__dfxtp_1
X_3396_ _2654_ _2906_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__and2_2
X_5135_ _0363_ _3040_ _3042_ _0366_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _2775_ _2716_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _2806_ _2735_ _0694_ _2739_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5968_ clknet_1_0__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__buf_1
X_4919_ _0407_ _3010_ BitStream_buffer.BS_buffer\[75\] _3013_ vssd1 vssd1 vccd1 vccd1
+ _1699_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5899_ _2474_ _2516_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6137__64 clknet_1_0__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__inv_2
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _2783_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__clkbuf_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _2714_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5822_ _2431_ _2445_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5753_ _2377_ _2310_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6045__141 clknet_1_1__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
X_4704_ BitStream_buffer.BS_buffer\[64\] _2980_ _2982_ BitStream_buffer.BS_buffer\[65\]
+ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5684_ exp_golomb_decoding.te_range\[2\] vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__inv_2
X_4635_ _2766_ _2616_ _2768_ _2623_ _1416_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _0464_ _2824_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__or2_1
X_6305_ net107 _0320_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3517_ BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__clkbuf_4
X_4497_ _2658_ _2998_ _0411_ _3001_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__o22ai_1
X_6236_ net38 _0251_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[31\] sky130_fd_sc_hd__dfxtp_2
X_3448_ _2680_ _2964_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__and2_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _2905_ _2909_ _2910_ _2912_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__o22ai_1
X_6167_ net129 _0182_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[109\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5118_ BitStream_buffer.BS_buffer\[58\] _2934_ BitStream_buffer.BS_buffer\[59\] _2937_
+ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__a221oi_1
X_5049_ _0398_ _3051_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4420_ _1161_ _1203_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6116__45 clknet_1_1__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__inv_2
XFILLER_0_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4351_ _2803_ BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__nand2_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4282_ _2996_ _2967_ _2999_ _2970_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__o22ai_1
X_6131__59 clknet_1_0__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__inv_2
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _2765_ _2766_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__nand2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__inv_2
X_3095_ net35 _2621_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5805_ _2427_ _2428_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__nand2_1
X_3997_ _0738_ _0784_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__nand3_1
X_5736_ _2360_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__inv_4
X_5667_ net8 BitStream_buffer.BS_buffer\[126\] _2266_ vssd1 vssd1 vccd1 vccd1 _2297_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4618_ _2910_ _0344_ _2914_ _0347_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5598_ _2249_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
X_4549_ _2737_ _2753_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6219_ net181 _0234_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[57\] sky130_fd_sc_hd__dfxtp_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3920_ _0445_ _2780_ _0706_ _0707_ _0708_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__o2111a_1
X_3851_ _0640_ _3026_ _0514_ _3030_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3782_ _2749_ BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__nand2_1
X_5521_ _2196_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5452_ _0404_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__clkbuf_2
X_5383_ _2102_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__nand2_2
X_4403_ _0358_ _3055_ _0660_ _3058_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__o22ai_1
X_4334_ _0694_ _2713_ _1116_ _1117_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o2111a_1
X_4265_ _0518_ _2876_ _3037_ _2879_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__a221oi_1
X_4196_ _0979_ _0980_ _0981_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__or4_1
X_3216_ _2749_ BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__nand2_1
X_3147_ _2680_ _2621_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__and2_2
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ _2610_ _2611_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5719_ _2315_ _2325_ _2312_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2593_ clknet_0__2593_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2593_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4050_ BitStream_buffer.BS_buffer\[122\] _2863_ BitStream_buffer.BS_buffer\[123\]
+ _2866_ _0837_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__a221oi_1
Xinput6 BitStream_buffer_input[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_4
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _0419_ _2655_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4883_ _2830_ BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__nand2_1
X_3903_ _2724_ _2714_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__nand2_1
X_3834_ BitStream_buffer.BS_buffer\[42\] _2949_ BitStream_buffer.BS_buffer\[43\] _2952_
+ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3765_ _0411_ _2646_ _0552_ _0553_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__o2111a_1
X_3696_ _0486_ _2909_ _2905_ _2912_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__o22ai_1
X_5504_ _2183_ _2171_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__and2_1
X_5435_ _2136_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5366_ _2089_ _2079_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__and2_1
X_4317_ _1102_ _0672_ _0674_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__a21oi_1
X_5297_ net14 BitStream_buffer.BS_buffer\[40\] _2024_ vssd1 vssd1 vccd1 vccd1 _2042_
+ sky130_fd_sc_hd__mux2_1
X_4248_ _2775_ _2797_ _1031_ _1032_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__o2111a_1
X_4179_ BitStream_buffer.BS_buffer\[59\] _2981_ _2983_ BitStream_buffer.BS_buffer\[60\]
+ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3550_ BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _1982_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_1
X_3481_ _3009_ _3011_ BitStream_buffer.BS_buffer\[63\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _3015_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _1922_ _1924_ _1926_ _1928_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__and4_1
X_4102_ _0880_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__nand2_1
X_5082_ _2786_ BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__nand2_1
X_4033_ _2803_ _2816_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4935_ _2914_ _0356_ _2917_ _0359_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_11 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _2760_ _2804_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3817_ _2892_ BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__nand2_1
X_4797_ _0492_ _2908_ _2939_ _2911_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__o22ai_1
X_3748_ _0366_ _0365_ BitStream_buffer.BS_buffer\[18\] _0369_ _0538_ vssd1 vssd1 vccd1
+ vccd1 _0539_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2595_ _2595_ vssd1 vssd1 vccd1 vccd1 clknet_0__2595_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3679_ _2856_ BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5418_ _2124_ _2079_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__and2_1
X_5349_ net14 BitStream_buffer.BS_buffer\[24\] _2061_ vssd1 vssd1 vccd1 vccd1 _2078_
+ sky130_fd_sc_hd__mux2_1
Xmax_cap35 _2628_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_2
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4720_ BitStream_buffer.BS_buffer\[19\] _0326_ _0328_ BitStream_buffer.BS_buffer\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__a22o_1
X_4651_ _2792_ _2728_ BitStream_buffer.BS_buffer\[105\] _2731_ _1432_ vssd1 vssd1
+ vccd1 vccd1 _1433_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3602_ _0333_ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__nand2_1
X_4582_ _2883_ _2896_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3533_ BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__buf_2
X_6252_ net54 _0267_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[47\] sky130_fd_sc_hd__dfxtp_2
X_3464_ _2997_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__buf_2
X_6183_ net145 _0198_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[93\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5203_ _1970_ _1952_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5134_ BitStream_buffer.BS_buffer\[18\] _3033_ _3035_ BitStream_buffer.BS_buffer\[19\]
+ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__a22o_1
X_3395_ _2928_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__buf_2
X_5065_ _1833_ _1837_ _1840_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4016_ _2733_ _2713_ _0801_ _0802_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__o2111a_1
X_5967_ clk vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__buf_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4918_ BitStream_buffer.BS_buffer\[68\] _2991_ BitStream_buffer.BS_buffer\[69\] _2994_
+ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _2421_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4849_ _2698_ _2645_ _1626_ _1627_ _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__o2111a_1
X_6022__120 clknet_1_1__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XFILLER_0_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__clkbuf_4
X_5821_ _2437_ _2444_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5752_ _2353_ _2327_ _2345_ _2608_ _2319_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__a311o_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4703_ _0632_ _2973_ _0505_ _2976_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__o22ai_1
X_5683_ net21 _2307_ net20 vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4634_ _2751_ _2629_ _0431_ _2636_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4565_ _2819_ _2838_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6304_ net106 _0319_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_3516_ _3049_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__buf_2
X_4496_ _1276_ _1277_ _1278_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__or4_1
X_6235_ net197 _0250_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc_previous\[6\] sky130_fd_sc_hd__dfxtp_2
X_3447_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__clkbuf_4
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__buf_4
X_6166_ net128 _0181_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[110\] sky130_fd_sc_hd__dfxtp_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _0632_ _2940_ _0505_ _2944_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__o22ai_1
X_5048_ _1795_ _1805_ _1826_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__nor3_1
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6029__126 clknet_1_0__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4350_ _2799_ BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nand2_1
X_3301_ _2834_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__buf_2
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ _1062_ _1064_ _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__nand3b_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__buf_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _2696_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__clkbuf_4
X_3094_ BitStream_buffer.pc\[2\] _2604_ _2627_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__nor3_2
XFILLER_0_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5804_ _2381_ BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1 vccd1
+ _2428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3996_ _0399_ _3044_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__nand2_1
X_5735_ _2341_ _2351_ _2346_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__nand3_4
XFILLER_0_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5666_ _2296_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4617_ _1394_ _1399_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5597_ _2248_ _2240_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__and2_1
X_4548_ _2749_ _2706_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nand2_1
X_4479_ _0727_ _2890_ _1260_ _1261_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__o2111a_1
X_6218_ net180 _0233_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[58\] sky130_fd_sc_hd__dfxtp_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ net111 _0164_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[127\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3850_ BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3781_ _2746_ _2766_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__nand2_1
X_5520_ _2194_ _2195_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5451_ net10 BitStream_buffer.BS_buffer\[60\] _2120_ vssd1 vssd1 vccd1 vccd1 _2147_
+ sky130_fd_sc_hd__mux2_1
X_5382_ BitStream_buffer.pc_previous\[3\] BitStream_buffer.exp_golomb_len\[3\] vssd1
+ vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__nand2_1
X_4402_ BitStream_buffer.BS_buffer\[19\] _3048_ _3050_ BitStream_buffer.BS_buffer\[20\]
+ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__a22o_1
X_4333_ _2724_ BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4264_ _0638_ _2882_ _0512_ _2885_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3215_ _2748_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4195_ _0521_ _0327_ _0329_ _3051_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__a22o_1
X_3146_ _2667_ _2619_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__nor2_4
X_3077_ _2607_ BitStream_buffer.pc_previous\[0\] vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__nand2_4
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5718_ BitStream_buffer.BitStream_buffer_output\[5\] _2342_ _1310_ _1414_ vssd1 vssd1
+ vccd1 vccd1 _2343_ sky130_fd_sc_hd__o211a_1
X_3979_ _0373_ _3055_ _0646_ _3058_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5649_ net19 vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__buf_2
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6058__152 clknet_1_1__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__2592_ clknet_0__2592_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2592_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 BitStream_buffer_input[15] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
X_4951_ _2649_ BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4882_ _2894_ _2812_ _1659_ _1660_ _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3902_ _2720_ BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__nand2_1
X_3833_ _0622_ _2955_ _0495_ _2959_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_52_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3764_ _2664_ _2661_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__or2_1
X_3695_ BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__inv_2
X_5503_ net10 BitStream_buffer.BS_buffer\[76\] _2156_ vssd1 vssd1 vccd1 vccd1 _2183_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5434_ _2135_ _2127_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5365_ net9 _0380_ _2060_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__mux2_1
X_4316_ BitStream_buffer.BitStream_buffer_output\[9\] vssd1 vssd1 vccd1 vccd1 _1102_
+ sky130_fd_sc_hd__inv_2
X_5296_ _2041_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__clkbuf_1
X_4247_ _2811_ _2808_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__or2_1
X_4178_ _0750_ _2974_ _0626_ _2977_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__o22ai_1
X_3129_ _2640_ _2646_ _2651_ _2657_ _2662_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3480_ _3013_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5150_ BitStream_buffer.BS_buffer\[42\] _0378_ BitStream_buffer.BS_buffer\[43\] _0382_
+ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__a221oi_1
X_4101_ _0882_ _0884_ _0886_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__and4_1
X_5081_ _2850_ _2783_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__or2_1
X_6086__18 clknet_1_1__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__inv_2
X_4032_ _2799_ _2820_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__nand2_1
X_5987__88 clknet_1_1__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
X_4934_ BitStream_buffer.BS_buffer\[36\] _0336_ BitStream_buffer.BS_buffer\[37\] _0340_
+ _1713_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _2733_ _2743_ _1642_ _1643_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3816_ _0400_ _2876_ BitStream_buffer.BS_buffer\[1\] _2879_ _0605_ vssd1 vssd1 vccd1
+ vccd1 _0606_ sky130_fd_sc_hd__a221oi_1
X_4796_ _1531_ _1546_ _1563_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3747_ _0537_ _0372_ _0370_ _0375_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2594_ _2594_ vssd1 vssd1 vccd1 vccd1 clknet_0__2594_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ _0468_ _2852_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5417_ net6 BitStream_buffer.BS_buffer\[49\] _2121_ vssd1 vssd1 vccd1 vccd1 _2124_
+ sky130_fd_sc_hd__mux2_1
X_5348_ _2077_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
X_5279_ _2029_ _1973_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap36 _2620_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
XFILLER_0_69_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4650_ _2811_ _2734_ _0459_ _2738_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__o22ai_1
X_3601_ _0349_ _0362_ _0377_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__and4_1
Xinput10 BitStream_buffer_input[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_4
X_4581_ _2892_ BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3532_ _3060_ _3062_ _3063_ _0323_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__o22ai_1
X_6251_ net53 _0266_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[16\] sky130_fd_sc_hd__dfxtp_1
X_3463_ net36 _2965_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__nand2_2
X_6182_ net144 _0197_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[94\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5202_ net13 _0325_ _1950_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__mux2_1
X_5133_ _0660_ _3025_ _0537_ _3029_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__o22ai_1
X_3394_ _2922_ _2643_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ _2736_ _2688_ BitStream_buffer.BS_buffer\[93\] _2692_ _1841_ vssd1 vssd1 vccd1
+ vccd1 _1842_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4015_ _2724_ _2736_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _2417_ _2574_ _2579_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5897_ _2514_ _2417_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__nand2_1
X_4917_ _0556_ _2997_ _0415_ _3000_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__o22ai_1
X_4848_ _0560_ _2660_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4779_ _2834_ BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5820_ _2403_ _2439_ _2443_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5751_ _2310_ _2375_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6006__105 clknet_1_0__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
X_4702_ _0508_ _2966_ _3009_ _2969_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5682_ _2306_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4633_ _2599_ _1413_ _1415_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4564_ _2815_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__nand2_1
X_6303_ net105 _0318_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3515_ _2695_ _3019_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__and2_2
X_6234_ net196 _0249_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc_previous\[5\] sky130_fd_sc_hd__dfxtp_1
X_4495_ BitStream_buffer.BS_buffer\[56\] _2986_ _2988_ BitStream_buffer.BS_buffer\[57\]
+ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__a22o_1
X_3446_ _2979_ _2677_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__nor2_2
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ net127 _0180_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[111\] sky130_fd_sc_hd__dfxtp_2
X_3377_ _2673_ _2907_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _1890_ _1891_ _1892_ _1893_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__or4_1
X_6052__147 clknet_1_1__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
X_5047_ _1816_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5949_ _2563_ _2564_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__nand2_1
XFILLER_0_47_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3300_ _2777_ _2687_ vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ BitStream_buffer.BS_buffer\[46\] _2949_ BitStream_buffer.BS_buffer\[47\] _2952_
+ _1065_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__a221oi_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _2764_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__buf_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _2695_ _2621_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__nand2_2
X_3093_ _2618_ _2626_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__nand2_4
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5803_ _2329_ _2360_ BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1
+ vccd1 _2427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3995_ _0749_ _0760_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__nor3_1
X_5734_ _2350_ _2358_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5665_ _2295_ _2285_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4616_ _1395_ _1396_ _1397_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5596_ net14 _2792_ _2230_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4547_ _2746_ _2714_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__nand2_1
X_4478_ _2850_ _2900_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__or2_1
X_3429_ BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__inv_2
X_6217_ net179 _0232_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[59\] sky130_fd_sc_hd__dfxtp_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ net110 _0163_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.buffer_index\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ clknet_1_1__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__buf_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6121__50 clknet_1_0__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__inv_2
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3780_ _2800_ _2729_ BitStream_buffer.BS_buffer\[97\] _2732_ _0569_ vssd1 vssd1 vccd1
+ vccd1 _0570_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5450_ _2146_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4401_ _1182_ _1183_ _1184_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5381_ BitStream_buffer.pc_previous\[3\] BitStream_buffer.exp_golomb_len\[3\] _2101_
+ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__o21ai_1
X_4332_ _2720_ BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__nand2_1
X_4263_ BitStream_buffer.BS_buffer\[124\] _2863_ BitStream_buffer.BS_buffer\[125\]
+ _2866_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6002_ clknet_1_0__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__buf_1
X_3214_ _2710_ _2643_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__nor2_2
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4194_ _0523_ _3062_ _3053_ _0323_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__o22ai_1
X_3145_ _2678_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3076_ _2608_ _2609_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ BitStream_buffer.BS_buffer\[15\] _3048_ _3050_ _0363_ vssd1 vssd1 vccd1 vccd1
+ _0767_ sky130_fd_sc_hd__a22o_1
X_5717_ BitStream_buffer.BitStream_buffer_output\[3\] BitStream_buffer.BitStream_buffer_output\[2\]
+ _1622_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5648_ net14 BitStream_buffer.BS_buffer\[120\] _2267_ vssd1 vssd1 vccd1 vccd1 _2284_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5579_ _2236_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__2591_ clknet_0__2591_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2591_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput8 BitStream_buffer_input[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_4
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4950_ _2756_ _2616_ _2725_ _2623_ _1728_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__a221oi_1
X_3901_ _0428_ _2717_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__or2_1
X_4881_ _2898_ _2823_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__or2_1
X_3832_ BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__inv_2
X_5502_ _2182_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__clkbuf_1
X_3763_ _2658_ _2656_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3694_ _0422_ _0443_ _0467_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5433_ net16 BitStream_buffer.BS_buffer\[54\] _2121_ vssd1 vssd1 vccd1 vccd1 _2135_
+ sky130_fd_sc_hd__mux2_1
X_5364_ _2088_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
X_4315_ _1057_ _1099_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__nand3_1
X_5295_ _2040_ _2034_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__and2_1
X_4246_ _2803_ _2792_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__nand2_1
X_6100__31 clknet_1_0__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__inv_2
X_4177_ _2999_ _2967_ _0858_ _2970_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__o22ai_1
X_3128_ _2658_ _2661_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4100_ BitStream_buffer.BS_buffer\[32\] _0379_ BitStream_buffer.BS_buffer\[33\] _0383_
+ _0887_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__a221oi_2
X_5080_ _1847_ _1849_ _1853_ _1857_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4031_ _2839_ _2780_ _0816_ _0817_ _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4933_ _0613_ _0343_ _0486_ _0346_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4864_ _0568_ _2752_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__or2_1
XANTENNA_13 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3815_ _0604_ _2882_ _0476_ _2885_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__o22ai_1
X_4795_ _1567_ _1569_ _1571_ _1575_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_24 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3746_ BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__inv_2
Xclkbuf_0__2593_ _2593_ vssd1 vssd1 vccd1 vccd1 clknet_0__2593_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3677_ BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
X_5416_ _2123_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
X_5347_ _2076_ _2055_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__and2_1
X_5278_ net5 BitStream_buffer.BS_buffer\[34\] _2024_ vssd1 vssd1 vccd1 vccd1 _2029_
+ sky130_fd_sc_hd__mux2_1
X_4229_ _0568_ _2713_ _1012_ _1013_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6091__22 clknet_1_1__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__inv_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3600_ BitStream_buffer.BS_buffer\[28\] _0379_ _0380_ _0383_ _0391_ vssd1 vssd1 vccd1
+ vccd1 _0392_ sky130_fd_sc_hd__a221oi_1
Xinput11 BitStream_buffer_input[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_4
X_4580_ BitStream_buffer.BS_buffer\[7\] _2876_ _0330_ _2879_ _1362_ vssd1 vssd1 vccd1
+ vccd1 _1363_ sky130_fd_sc_hd__a221oi_1
X_5992__92 clknet_1_0__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
XFILLER_0_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3531_ _0322_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6250_ net52 _0265_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[17\] sky130_fd_sc_hd__dfxtp_1
X_3462_ BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__inv_2
X_3393_ BitStream_buffer.BS_buffer\[38\] _2924_ _2926_ BitStream_buffer.BS_buffer\[39\]
+ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__a22o_1
X_5201_ _1969_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
X_6181_ net143 _0196_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[95\] sky130_fd_sc_hd__dfxtp_2
X_5132_ _3053_ _3021_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5063_ _2715_ _2696_ _0423_ _2701_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6075__8 clknet_1_1__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__inv_2
X_4014_ _2720_ BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5965_ net18 _2310_ _2606_ _2567_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5896_ _2512_ _2513_ _2375_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__o21ai_1
X_4916_ _1692_ _1693_ _1694_ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4847_ _2694_ _2655_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4778_ _2830_ BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__nand2_1
X_3729_ _0513_ _0515_ _0517_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6128__56 clknet_1_0__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__inv_2
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5750_ _2374_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5681_ net18 net17 vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4701_ _1478_ _1480_ _1482_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4632_ _1414_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4563_ _0445_ _2797_ _1343_ _1344_ _1345_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__o2111a_1
X_6302_ net104 _0317_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3514_ _3047_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__buf_2
X_4494_ BitStream_buffer.BS_buffer\[62\] _2981_ _2983_ BitStream_buffer.BS_buffer\[63\]
+ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__a22o_1
X_6233_ net195 _0248_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc_previous\[4\] sky130_fd_sc_hd__dfxtp_2
X_3445_ _2964_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__inv_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__inv_2
X_6164_ net126 _0179_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[112\] sky130_fd_sc_hd__dfxtp_2
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ BitStream_buffer.BS_buffer\[46\] _2928_ _2930_ BitStream_buffer.BS_buffer\[47\]
+ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__a22o_1
X_5046_ _1818_ _1820_ _1822_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5948_ _2529_ _2516_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5879_ _2492_ _2496_ _2371_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__nand3_1
XFILLER_0_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5971__73 clknet_1_1__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__inv_2
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _2710_ _2672_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__nor2_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _2685_ _2627_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nor2_4
X_3092_ BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__inv_2
X_5802_ _2422_ _2425_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3994_ _0773_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5733_ BitStream_buffer.BitStream_buffer_output\[7\] _2354_ _2357_ vssd1 vssd1 vccd1
+ vccd1 _2358_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5664_ net9 BitStream_buffer.BS_buffer\[125\] _2266_ vssd1 vssd1 vccd1 vccd1 _2295_
+ sky130_fd_sc_hd__mux2_1
X_4615_ BitStream_buffer.BS_buffer\[18\] _0327_ _0329_ _0366_ vssd1 vssd1 vccd1 vccd1
+ _1398_ sky130_fd_sc_hd__a22o_1
X_5595_ _2247_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
X_4546_ BitStream_buffer.BS_buffer\[103\] _2729_ _2792_ _2732_ _1328_ vssd1 vssd1
+ vccd1 vccd1 _1329_ sky130_fd_sc_hd__a221oi_1
X_6107__37 clknet_1_1__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__inv_2
X_4477_ _2845_ _2896_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__or2_1
X_3428_ _2933_ _2947_ _2961_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__nand3b_1
X_6216_ net178 _0231_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[60\] sky130_fd_sc_hd__dfxtp_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ net109 _0162_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.buffer_index\[5\] sky130_fd_sc_hd__dfxtp_1
X_3359_ _2892_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__nand2_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5029_ _0366_ _3033_ _3035_ BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1
+ _1808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4400_ _0325_ _3041_ _3043_ _0527_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5380_ _2098_ _2099_ _2100_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4331_ _0453_ _2717_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__or2_1
X_4262_ _2845_ _2869_ _0468_ _2872_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3213_ _2746_ BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4193_ _0537_ _3055_ _0370_ _3058_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__o22ai_1
X_3144_ _2603_ _2677_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__nor2_2
X_3075_ BitStream_buffer.pc_previous\[0\] vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3977_ _0762_ _0763_ _0764_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5716_ _2340_ _2311_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5647_ _2283_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
X_5578_ _2235_ _2216_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__and2_1
X_4529_ _0431_ _2630_ _2742_ _2637_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__o22ai_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__2590_ clknet_0__2590_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2590_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 BitStream_buffer_input[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_4
XFILLER_0_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4880_ _2818_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__nand2_1
X_3900_ _0678_ _0682_ _0685_ _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__and4_1
X_3831_ BitStream_buffer.BS_buffer\[46\] _2935_ BitStream_buffer.BS_buffer\[47\] _2938_
+ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3762_ _2650_ BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5501_ _2181_ _2171_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3693_ _0472_ _0475_ _0478_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5432_ _2134_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
X_5363_ _2087_ _2079_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _0399_ _0516_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nand2_1
X_5294_ net15 BitStream_buffer.BS_buffer\[39\] _2024_ vssd1 vssd1 vccd1 vccd1 _2040_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4245_ _2799_ _2816_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__nand2_1
X_4176_ _0958_ _0960_ _0962_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__nand3b_1
X_3127_ _2660_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4030_ _2791_ _2832_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4932_ _1706_ _1711_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4863_ _2748_ _2736_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__nand2_1
XANTENNA_14 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4794_ _2845_ _2889_ _1572_ _1573_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__o2111a_1
X_3814_ BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__inv_2
XANTENNA_25 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ BitStream_buffer.BS_buffer\[21\] _0351_ BitStream_buffer.BS_buffer\[22\] _0354_
+ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2592_ _2592_ vssd1 vssd1 vccd1 vccd1 clknet_0__2592_ sky130_fd_sc_hd__clkbuf_16
X_5415_ _2122_ _2079_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__and2_1
X_3676_ _0449_ _0455_ _0461_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5346_ net15 BitStream_buffer.BS_buffer\[23\] _2061_ vssd1 vssd1 vccd1 vccd1 _2076_
+ sky130_fd_sc_hd__mux2_1
X_5277_ _2028_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
X_4228_ _2724_ BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__nand2_1
X_4159_ _0512_ _2882_ _3018_ _2885_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput12 BitStream_buffer_input[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_8
X_3530_ _2957_ _3020_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__nand2_2
X_3461_ _2994_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__buf_2
X_5200_ _1968_ _1952_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__and2_1
X_3392_ _2925_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__clkbuf_4
X_6180_ net142 _0195_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[96\] sky130_fd_sc_hd__dfxtp_1
X_5131_ _1904_ _1906_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__nand3b_1
X_5062_ _1838_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4013_ _0568_ _2717_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5964_ _2577_ _2578_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__nand2_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5895_ _2511_ _2504_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__and2_1
X_4915_ BitStream_buffer.BS_buffer\[60\] _2985_ _2987_ BitStream_buffer.BS_buffer\[61\]
+ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4846_ _2649_ BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4777_ _0481_ _2812_ _1555_ _1556_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3728_ _3044_ _3041_ _3043_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__a22o_1
X_3659_ _2820_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
X_5329_ _2064_ _2055_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5680_ _2305_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_4700_ BitStream_buffer.BS_buffer\[50\] _2948_ BitStream_buffer.BS_buffer\[51\] _2951_
+ _1481_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4631_ BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1 vccd1 _1414_
+ sky130_fd_sc_hd__inv_2
X_4562_ _0444_ _2808_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__or2_1
X_6301_ net103 _0316_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3513_ _3032_ _2699_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__nor2_2
X_4493_ _2996_ _2974_ _2999_ _2977_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__o22ai_1
X_6232_ net194 _0247_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc_previous\[3\] sky130_fd_sc_hd__dfxtp_1
X_3444_ _2972_ _2974_ _2975_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__o22ai_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ net125 _0178_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[113\] sky130_fd_sc_hd__dfxtp_2
X_3375_ _2908_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__clkbuf_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ BitStream_buffer.BS_buffer\[52\] _2923_ _2925_ BitStream_buffer.BS_buffer\[53\]
+ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__a22o_1
X_5045_ BitStream_buffer.BS_buffer\[41\] _0378_ BitStream_buffer.BS_buffer\[42\] _0382_
+ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5947_ _2554_ _2417_ _2562_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5878_ _2494_ _2495_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__nand2_1
X_4829_ BitStream_buffer.BS_buffer\[35\] _0336_ BitStream_buffer.BS_buffer\[36\] _0340_
+ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__inv_2
Xhold1 net30 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__inv_2
X_6012__111 clknet_1_1__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5801_ _2423_ _2424_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5732_ _2356_ _2353_ _0894_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__nand3_1
X_3993_ _0775_ _0777_ _0779_ _0781_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ _2294_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4614_ _0537_ _3062_ _0370_ _0323_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__o22ai_1
X_5594_ _2246_ _2240_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__and2_1
X_4545_ _0459_ _2735_ _2822_ _2739_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__o22ai_1
X_4476_ _2892_ BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nand2_1
X_6215_ net177 _0230_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[61\] sky130_fd_sc_hd__dfxtp_2
X_3427_ BitStream_buffer.BS_buffer\[40\] _2949_ BitStream_buffer.BS_buffer\[41\] _2952_
+ _2960_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__a221oi_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ net108 _0161_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.buffer_index\[4\] sky130_fd_sc_hd__dfxtp_1
X_3358_ _2891_ vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__buf_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3289_ _2668_ _2778_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__nand2_1
X_5028_ _0537_ _3025_ _0370_ _3029_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ _1105_ _1109_ _1112_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__and4_1
X_4261_ _3018_ _2849_ _1044_ _1045_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3212_ _2745_ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4192_ _0366_ _3048_ _3050_ BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1
+ _0979_ sky130_fd_sc_hd__a22o_1
X_3143_ _2647_ _2666_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__nand2_4
X_3074_ _2607_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3976_ _3037_ _3041_ _3043_ _0516_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__a22o_1
X_5715_ _2338_ _2339_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5646_ _2282_ _2261_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5577_ net5 _2804_ _2230_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__mux2_1
X_4528_ _2599_ _1309_ _1311_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__o21a_1
X_6019__117 clknet_1_1__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
X_4459_ _2815_ _2836_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__nand2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065__159 clknet_1_0__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6098__29 clknet_1_0__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__inv_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5999__99 clknet_1_1__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3830_ _0619_ _2941_ _0492_ _2945_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__o22ai_1
X_3761_ BitStream_buffer.BS_buffer\[76\] _2617_ BitStream_buffer.BS_buffer\[77\] _2624_
+ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5500_ net11 BitStream_buffer.BS_buffer\[75\] _2156_ vssd1 vssd1 vccd1 vccd1 _2181_
+ sky130_fd_sc_hd__mux2_1
X_3692_ _2898_ _2890_ _0479_ _0480_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__o2111a_1
X_5431_ _2133_ _2127_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__and2_1
X_5362_ net10 BitStream_buffer.BS_buffer\[28\] _2060_ vssd1 vssd1 vccd1 vccd1 _2087_
+ sky130_fd_sc_hd__mux2_1
X_4313_ _1067_ _1077_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__nor3_1
X_5293_ _2039_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
X_4244_ _2827_ _2780_ _1027_ _1028_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__o2111a_1
X_4175_ BitStream_buffer.BS_buffer\[45\] _2949_ BitStream_buffer.BS_buffer\[46\] _2952_
+ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__a221oi_1
X_3126_ _2659_ _2621_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__nand2_1
X_3959_ BitStream_buffer.BS_buffer\[43\] _2949_ BitStream_buffer.BS_buffer\[44\] _2952_
+ _0747_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5629_ _2271_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5980_ clknet_1_0__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__buf_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4931_ _1707_ _1708_ _1709_ _1710_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__or4_1
X_6048__143 clknet_1_0__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
X_4862_ _2745_ BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__nand2_1
X_3813_ BitStream_buffer.BS_buffer\[120\] _2863_ BitStream_buffer.BS_buffer\[121\]
+ _2866_ _0602_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__a221oi_1
X_4793_ _2883_ _2899_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__or2_1
XANTENNA_15 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__2591_ _2591_ vssd1 vssd1 vccd1 vccd1 clknet_0__2591_ sky130_fd_sc_hd__clkbuf_16
X_3744_ _0534_ _0357_ _0355_ _0360_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3675_ _2888_ _2829_ _0462_ _0463_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__o2111a_1
X_5414_ net7 BitStream_buffer.BS_buffer\[48\] _2121_ vssd1 vssd1 vccd1 vccd1 _2122_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5345_ _2075_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5276_ _2027_ _1973_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__and2_1
X_4227_ _2720_ _2800_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nand2_1
X_4158_ BitStream_buffer.BS_buffer\[123\] _2863_ BitStream_buffer.BS_buffer\[124\]
+ _2866_ _0944_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__a221oi_1
X_4089_ _3053_ _3062_ _3056_ _0323_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__o22ai_1
X_3109_ _2641_ _2642_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__nand2_4
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 BitStream_buffer_input[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_4
XFILLER_0_12_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3460_ _2993_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__clkbuf_2
X_3391_ _2680_ _2906_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__and2_2
X_5130_ BitStream_buffer.BS_buffer\[74\] _3004_ BitStream_buffer.BS_buffer\[75\] _3007_
+ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__a221oi_1
X_5061_ _2766_ _2678_ _2681_ _2768_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__a22o_1
X_4012_ _0790_ _0794_ _0797_ _0799_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5963_ net18 _2310_ _2606_ _2556_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4914_ BitStream_buffer.BS_buffer\[66\] _2980_ _2982_ BitStream_buffer.BS_buffer\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5894_ _2504_ _2511_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4845_ _2762_ _2616_ _2756_ _2623_ _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4776_ _2888_ _2823_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3727_ BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3658_ _0444_ _2780_ _0446_ _0447_ _0448_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__o2111a_1
X_3589_ _2695_ _0334_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__and2_1
X_5328_ net6 _0366_ _2061_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__mux2_1
X_5259_ net33 _2012_ _2014_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4630_ _1369_ _1411_ _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6300_ net102 _0315_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BitStream_buffer_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_4561_ _2803_ _2781_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3512_ _3023_ _3031_ _3038_ _3045_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__or4_1
X_4492_ _0632_ _2967_ _0505_ _2970_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__o22ai_1
X_6231_ net193 _0246_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc_previous\[2\] sky130_fd_sc_hd__dfxtp_1
X_3443_ _2976_ vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__buf_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ net124 _0177_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[114\] sky130_fd_sc_hd__dfxtp_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3374_ _2668_ _2907_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__nand2_2
X_5113_ _0619_ _2915_ _0492_ _2919_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__o22ai_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _0495_ _0385_ _2953_ _0389_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5946_ _2561_ _2374_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__nand2_1
X_5877_ _2491_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4828_ _0486_ _0343_ _2905_ _0346_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4759_ _0428_ _2752_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__or2_1
X_6133__61 clknet_1_0__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__inv_2
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 _1942_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _2623_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__clkbuf_4
X_5800_ _2361_ _1726_ _2328_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__nand3_1
X_3992_ BitStream_buffer.BS_buffer\[32\] _0382_ BitStream_buffer.BS_buffer\[31\] _0379_
+ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__a221oi_1
X_5731_ _2355_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2597_ clknet_0__2597_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2597_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5662_ _2293_ _2285_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4613_ _0534_ _3055_ _0355_ _3058_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__o22ai_1
X_5593_ net15 BitStream_buffer.BS_buffer\[103\] _2230_ vssd1 vssd1 vccd1 vccd1 _2246_
+ sky130_fd_sc_hd__mux2_1
X_4544_ _0453_ _2713_ _1324_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__o2111a_1
X_6214_ net176 _0229_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[62\] sky130_fd_sc_hd__dfxtp_2
X_4475_ _0516_ _2876_ BitStream_buffer.BS_buffer\[7\] _2879_ _1258_ vssd1 vssd1 vccd1
+ vccd1 _1259_ sky130_fd_sc_hd__a221oi_1
X_3426_ _2953_ _2955_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__o22ai_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _2854_ _2648_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__nor2_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _3056_ _3021_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__nor2_1
X_3288_ BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5929_ _2542_ _2544_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6042__138 clknet_1_1__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4260_ _2859_ BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nand2_1
X_4191_ _0974_ _0975_ _0976_ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__or4_1
X_3211_ _2710_ _2648_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__nor2_2
X_3142_ _2664_ _2670_ _2671_ _2675_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__o22ai_1
X_3073_ _2605_ _2606_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__nand2_4
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3975_ BitStream_buffer.BS_buffer\[7\] _3034_ _3036_ _0330_ vssd1 vssd1 vccd1 vccd1
+ _0764_ sky130_fd_sc_hd__a22o_1
X_5714_ _0787_ BitStream_buffer.BitStream_buffer_output\[11\] BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5645_ net15 BitStream_buffer.BS_buffer\[119\] _2267_ vssd1 vssd1 vccd1 vccd1 _2282_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5576_ _2234_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4527_ _1310_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4458_ _2782_ _2797_ _1239_ _1240_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__o2111a_1
X_3409_ _2687_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__inv_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ BitStream_buffer.BS_buffer\[61\] _2981_ _2983_ BitStream_buffer.BS_buffer\[62\]
+ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__a22o_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3760_ _0549_ _2630_ _0407_ _2637_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3691_ _0481_ _2900_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5430_ net2 BitStream_buffer.BS_buffer\[53\] _2121_ vssd1 vssd1 vccd1 vccd1 _2133_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _2086_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _2038_ _2034_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__and2_1
X_4312_ _1088_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nand2_1
X_4243_ _2791_ _2836_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nand2_1
X_4174_ _0492_ _2955_ _2939_ _2959_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__o22ai_1
X_3125_ _2653_ _2619_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__nor2_4
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6025__122 clknet_1_1__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
X_3958_ _2942_ _2955_ _0622_ _2959_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3889_ BitStream_buffer.BS_buffer\[77\] _2617_ BitStream_buffer.BS_buffer\[78\] _2624_
+ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__a221oi_1
X_5628_ _2270_ _2261_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5559_ net9 BitStream_buffer.BS_buffer\[93\] _2192_ vssd1 vssd1 vccd1 vccd1 _2222_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4930_ BitStream_buffer.BS_buffer\[21\] _0326_ _0328_ BitStream_buffer.BS_buffer\[20\]
+ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4861_ _2788_ _2728_ _2781_ _2731_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3812_ _0601_ _2869_ _0473_ _2872_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4792_ _0476_ _2895_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__or2_1
XANTENNA_16 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2590_ _2590_ vssd1 vssd1 vccd1 vccd1 clknet_0__2590_ sky130_fd_sc_hd__clkbuf_16
X_3743_ BitStream_buffer.BS_buffer\[24\] vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3674_ _0464_ _2841_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5413_ _2120_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__buf_4
X_5344_ _2074_ _2055_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__and2_1
X_5275_ net6 BitStream_buffer.BS_buffer\[33\] _2024_ vssd1 vssd1 vccd1 vccd1 _2027_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4226_ _2806_ _2717_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__or2_1
X_4157_ _0468_ _2869_ _2850_ _2872_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__o22ai_1
X_3108_ BitStream_buffer.pc\[2\] BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1
+ _2642_ sky130_fd_sc_hd__nor2_2
XFILLER_0_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4088_ _0370_ _3055_ _0373_ _3058_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 BitStream_buffer_input[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3390_ _2923_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__clkbuf_4
X_5060_ _2751_ _2669_ _0431_ _2674_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__o22ai_1
X_4011_ BitStream_buffer.BS_buffer\[82\] _2689_ BitStream_buffer.BS_buffer\[83\] _2693_
+ _0798_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6082__14 clknet_1_0__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__inv_2
XFILLER_0_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5962_ _2576_ _2417_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__nand2_1
X_4913_ _0508_ _2973_ _3009_ _2976_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__o22ai_1
X_5893_ _2472_ _2510_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4844_ _2769_ _2629_ _0434_ _2636_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5983__84 clknet_1_0__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__inv_2
X_4775_ _2818_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__nand2_1
X_3726_ BitStream_buffer.BS_buffer\[5\] _3034_ _3036_ _0516_ vssd1 vssd1 vccd1 vccd1
+ _0517_ sky130_fd_sc_hd__a22o_1
X_3657_ _2791_ BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__nand2_1
X_3588_ BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__clkbuf_4
X_5327_ _2063_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
X_5258_ _0675_ _2014_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__nor2_1
X_5189_ _1961_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
X_4209_ _0399_ _3037_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4560_ _2799_ BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6119__48 clknet_1_0__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__inv_2
XFILLER_0_12_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3511_ _3039_ _3041_ _3043_ _3044_ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__a22o_1
X_4491_ _1270_ _1272_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand3b_1
X_6230_ net192 _0245_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc_previous\[1\] sky130_fd_sc_hd__dfxtp_1
X_3442_ _2918_ _2965_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__nand2_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ net123 _0176_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[115\] sky130_fd_sc_hd__dfxtp_2
X_3373_ _2906_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__clkbuf_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _2972_ _2908_ _2975_ _2911_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__o22ai_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5043_ _0380_ _0364_ _0387_ _0368_ _1821_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5945_ _2558_ _2560_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5876_ _2493_ _2453_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4827_ _1602_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4758_ _2748_ _2714_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__nand2_1
X_4689_ _0468_ _2889_ _1468_ _1469_ _1470_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3709_ _0499_ _2967_ _2963_ _2970_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 _1943_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3991_ _2917_ _0386_ _0663_ _0390_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5730_ _2351_ _2326_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2596_ clknet_0__2596_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2596_
+ sky130_fd_sc_hd__clkbuf_16
X_5661_ net10 BitStream_buffer.BS_buffer\[124\] _2266_ vssd1 vssd1 vccd1 vccd1 _2293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4612_ BitStream_buffer.BS_buffer\[21\] _3048_ _3050_ BitStream_buffer.BS_buffer\[22\]
+ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__a22o_1
X_5592_ _2245_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4543_ _2724_ BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__nand2_1
X_4474_ _0869_ _2882_ _0761_ _2885_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__o22ai_1
X_6213_ net175 _0228_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[63\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3425_ _2958_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__clkbuf_4
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _2889_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__buf_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _2819_ _2820_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__nand2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5026_ _1800_ _1802_ _1804_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__nand3b_1
X_5928_ _2543_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5859_ _2480_ vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ BitStream_buffer.BS_buffer\[7\] _3041_ _3043_ _0330_ vssd1 vssd1 vccd1 vccd1
+ _0977_ sky130_fd_sc_hd__a22o_1
X_3210_ _2743_ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__buf_2
X_3141_ _2674_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__clkbuf_4
X_3072_ net17 vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3974_ _3063_ _3026_ _0640_ _3030_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_72_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5713_ _2337_ _2316_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5644_ _2281_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5575_ _2233_ _2216_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__and2_1
X_4526_ BitStream_buffer.BitStream_buffer_output\[7\] vssd1 vssd1 vccd1 vccd1 _1310_
+ sky130_fd_sc_hd__inv_2
X_4457_ _2775_ _2808_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__or2_1
X_3408_ BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__inv_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4388_ _2999_ _2974_ _0858_ _2977_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__o22ai_1
X_3339_ _2867_ _2869_ _2870_ _2872_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__o22ai_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ BitStream_buffer.BS_buffer\[51\] _2923_ _2925_ BitStream_buffer.BS_buffer\[52\]
+ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3690_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5360_ _2085_ _2079_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__and2_1
X_4311_ _1090_ _1092_ _1094_ _1096_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__and4_1
X_5291_ net16 BitStream_buffer.BS_buffer\[38\] _2024_ vssd1 vssd1 vccd1 vccd1 _2038_
+ sky130_fd_sc_hd__mux2_1
X_4242_ _2787_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nand2_1
X_4173_ BitStream_buffer.BS_buffer\[49\] _2935_ BitStream_buffer.BS_buffer\[50\] _2938_
+ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__a221oi_2
X_3124_ BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3957_ BitStream_buffer.BS_buffer\[47\] _2935_ BitStream_buffer.BS_buffer\[48\] _2938_
+ _0745_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3888_ _2698_ _2630_ _0549_ _2637_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__o22ai_1
X_5627_ net6 BitStream_buffer.BS_buffer\[113\] _2267_ vssd1 vssd1 vccd1 vccd1 _2270_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5558_ _2221_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4509_ _0370_ _3062_ _0373_ _0323_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5489_ _2173_ _2171_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__and2_1
X_6088__20 clknet_1_1__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__inv_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989__90 clknet_1_1__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4860_ _2775_ _2734_ _0456_ _2738_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__o22ai_1
X_3811_ BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__inv_2
XANTENNA_28 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4791_ _2891_ BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3742_ BitStream_buffer.BS_buffer\[25\] _0337_ BitStream_buffer.BS_buffer\[26\] _0341_
+ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3673_ _2836_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
X_5412_ _2119_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5343_ net16 BitStream_buffer.BS_buffer\[22\] _2061_ vssd1 vssd1 vccd1 vccd1 _2074_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5274_ _2026_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
X_4225_ _1001_ _1005_ _1008_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__and4_1
X_4156_ _0730_ _2849_ _0940_ _0941_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__o2111a_1
X_3107_ _2632_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__inv_2
X_4087_ _0363_ _3048_ _3050_ _0366_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4989_ _2834_ BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 BitStream_buffer_input[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4010_ _2742_ _2697_ _0686_ _2702_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__o22ai_1
X_5961_ _2571_ _2575_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__nand2_1
X_4912_ _2652_ _2966_ _2640_ _2969_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__o22ai_1
X_5892_ _2416_ _2447_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__nor2_1
X_4843_ _0672_ _1621_ _1623_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4774_ _2814_ BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nand2_1
X_3725_ BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3656_ _2787_ _2781_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3587_ _0378_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5326_ _2062_ _2055_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__and2_1
X_5257_ _2013_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__inv_2
X_4208_ _0963_ _0973_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__nor3_1
X_5188_ _1960_ _1952_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__and2_1
X_4139_ _0464_ _2780_ _0923_ _0924_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3510_ BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4490_ BitStream_buffer.BS_buffer\[48\] _2949_ BitStream_buffer.BS_buffer\[49\] _2952_
+ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__a221oi_1
X_3441_ BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__inv_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ net122 _0175_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[116\] sky130_fd_sc_hd__dfxtp_2
X_3372_ _2708_ _2600_ BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__and3_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5111_ _1843_ _1858_ _1875_ _1888_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__and4_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _0540_ _0371_ _0384_ _0374_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5944_ _2508_ _2559_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__nand2_1
X_5875_ _2429_ _2455_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _1603_ _1604_ _1605_ _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4757_ _2745_ BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4688_ _2845_ _2899_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3708_ BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__inv_2
X_3639_ BitStream_buffer.BS_buffer\[95\] _2729_ _2800_ _2732_ _0429_ vssd1 vssd1 vccd1
+ vccd1 _0430_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ net10 BitStream_buffer.BS_buffer\[44\] _2023_ vssd1 vssd1 vccd1 vccd1 _2050_
+ sky130_fd_sc_hd__mux2_1
X_6289_ net91 _0304_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124__52 clknet_1_1__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__inv_2
Xhold4 _1944_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3990_ BitStream_buffer.BS_buffer\[19\] _0365_ BitStream_buffer.BS_buffer\[20\] _0369_
+ _0778_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _2292_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2595_ clknet_0__2595_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2595_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4611_ _1390_ _1391_ _1392_ _1393_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5591_ _2244_ _2240_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4542_ _2720_ BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nand2_1
X_4473_ BitStream_buffer.BS_buffer\[126\] _2863_ BitStream_buffer.BS_buffer\[127\]
+ _2866_ _1256_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__a221oi_1
X_3424_ _2957_ _2907_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6212_ net174 _0227_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[64\] sky130_fd_sc_hd__dfxtp_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3355_ _2644_ _2847_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__nand2_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3286_ BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__clkbuf_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ BitStream_buffer.BS_buffer\[73\] _3004_ BitStream_buffer.BS_buffer\[74\] _3007_
+ _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5927_ _1310_ _2366_ _1102_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ net20 net21 vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__nand2_1
X_5789_ _2392_ _2413_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__nand2_1
X_4809_ BitStream_buffer.BS_buffer\[65\] _2980_ _2982_ BitStream_buffer.BS_buffer\[66\]
+ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3140_ _2673_ _2621_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__nand2_2
X_3071_ net18 vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _2336_ _1102_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__nand2_1
X_3973_ _0761_ _3022_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5643_ _2280_ _2261_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5574_ net6 BitStream_buffer.BS_buffer\[97\] _2230_ vssd1 vssd1 vccd1 vccd1 _2233_
+ sky130_fd_sc_hd__mux2_1
X_4525_ _1265_ _1307_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nand3_1
X_4456_ _2803_ _2788_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__nand2_1
X_3407_ _2940_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__buf_2
X_4387_ _0505_ _2967_ _2996_ _2970_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__o22ai_1
X_6103__33 clknet_1_1__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__inv_2
X_3338_ _2871_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__buf_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ clknet_1_1__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__buf_1
X_3269_ _2802_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__clkbuf_4
X_5008_ _0492_ _2915_ _2939_ _2919_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5290_ _2037_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__clkbuf_1
X_4310_ BitStream_buffer.BS_buffer\[34\] _0379_ BitStream_buffer.BS_buffer\[35\] _0383_
+ _1095_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _2898_ _2784_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__or2_1
X_4172_ _2968_ _2941_ _2972_ _2945_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__o22ai_1
X_3123_ _2652_ _2656_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__or2_1
X_3956_ _2975_ _2941_ _0619_ _2945_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3887_ _2599_ _0670_ _0676_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__o21a_1
X_5626_ _2269_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5557_ _2220_ _2216_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__and2_1
X_5488_ net15 BitStream_buffer.BS_buffer\[71\] _2157_ vssd1 vssd1 vccd1 vccd1 _2173_
+ sky130_fd_sc_hd__mux2_1
X_4508_ _0355_ _3055_ _0358_ _3058_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__o22ai_1
X_4439_ _2806_ _2713_ _1220_ _1221_ _1222_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6009__108 clknet_1_1__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
X_3810_ _2880_ _2849_ _0597_ _0598_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4790_ _0325_ _2875_ _0527_ _2878_ _1570_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3741_ _0531_ _0344_ _0342_ _0347_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__o22ai_1
XANTENNA_18 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3672_ _2835_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__nand2_1
X_5411_ BitStream_buffer.buffer_index\[6\] _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__or2_1
X_5342_ _2073_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5273_ _2025_ _1973_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__and2_1
X_4224_ _2766_ _2689_ _2768_ _2693_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__a221oi_1
X_4155_ _2859_ BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__nand2_1
X_3106_ BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__inv_2
X_4086_ _0870_ _0871_ _0872_ _0873_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4988_ _2830_ BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3939_ _0727_ _2869_ _0601_ _2872_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5609_ _2256_ _2240_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 BitStream_buffer_input[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_4
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5960_ _2573_ _2574_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__nand2_1
X_5891_ _2506_ _2508_ _2374_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__o21a_1
X_4911_ _1686_ _1688_ _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4842_ _1622_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _0464_ _2796_ _1551_ _1552_ _1553_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o2111a_1
X_3724_ _0514_ _3026_ _3024_ _3030_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__o22ai_1
X_3655_ _0445_ _2784_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3586_ _0335_ _2699_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5325_ net7 _0363_ _2061_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__mux2_1
X_5256_ _2012_ net33 net34 vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ _0984_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5187_ net3 _0518_ _1950_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__mux2_1
X_4138_ _2791_ _2838_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__nand2_1
X_4069_ _0852_ _0854_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6038__134 clknet_1_0__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3440_ _2973_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__clkbuf_4
X_3371_ BitStream_buffer.BS_buffer\[37\] vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__inv_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ clknet_1_1__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__buf_1
XFILLER_0_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5110_ _1879_ _1881_ _1883_ _1887_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__and4_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ BitStream_buffer.BS_buffer\[33\] _0350_ BitStream_buffer.BS_buffer\[34\] _0353_
+ _1819_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5943_ _2548_ _2529_ _2415_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__o21ai_1
X_5874_ _2489_ _2491_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__nand2_1
X_4825_ BitStream_buffer.BS_buffer\[20\] _0326_ _0328_ BitStream_buffer.BS_buffer\[19\]
+ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4756_ BitStream_buffer.BS_buffer\[105\] _2728_ _2788_ _2731_ _1536_ vssd1 vssd1
+ vccd1 vccd1 _1537_ sky130_fd_sc_hd__a221oi_1
X_4687_ _2880_ _2895_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__or2_1
X_3707_ _0491_ _0494_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3638_ _0428_ _2735_ _2733_ _2739_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__o22ai_1
X_3569_ _0355_ _0357_ _0358_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__o22ai_1
X_5308_ _2049_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__clkbuf_1
X_6288_ net90 _0303_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[3\] sky130_fd_sc_hd__dfxtp_1
X_5239_ net28 _1941_ _1942_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2594_ clknet_0__2594_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2594_
+ sky130_fd_sc_hd__clkbuf_16
X_4610_ _0650_ _3041_ _3043_ _0770_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5590_ net16 _2816_ _2230_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__mux2_1
X_4541_ _0450_ _2717_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4472_ _2880_ _2869_ _2883_ _2872_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6211_ net173 _0226_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[65\] sky130_fd_sc_hd__dfxtp_2
X_3423_ _2615_ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__inv_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__inv_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _2818_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__clkbuf_4
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _0549_ _3010_ BitStream_buffer.BS_buffer\[76\] _3013_ vssd1 vssd1 vccd1 vccd1
+ _1803_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5926_ _2489_ _2541_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5857_ _2478_ _2479_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__nand2_1
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5788_ _2401_ _2412_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__nor2_1
X_4808_ _3009_ _2973_ _0632_ _2976_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4739_ _0434_ _2629_ _2751_ _2636_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3070_ BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5711_ _2335_ _1206_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__nand2_1
X_3972_ BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5642_ net16 BitStream_buffer.BS_buffer\[118\] _2267_ vssd1 vssd1 vccd1 vccd1 _2280_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5573_ _2232_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4524_ _0399_ _0330_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4455_ _2799_ _2792_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__nand2_1
X_4386_ _1166_ _1168_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nand3b_1
X_3406_ _2690_ _2907_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3337_ _2673_ _2847_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__nand2_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _2777_ _2648_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__nor2_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _2975_ _2908_ _0619_ _2911_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__o22ai_1
X_3199_ BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5909_ _2524_ _2525_ _2371_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4240_ _1015_ _1017_ _1021_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__and4_1
X_4171_ _0954_ _0955_ _0956_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__or4_1
X_3122_ _2655_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ _0740_ _0741_ _0742_ _0743_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3886_ _0671_ _0672_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__a21oi_1
X_5625_ _2268_ _2261_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5556_ net10 _2736_ _2192_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__mux2_1
X_5487_ _2172_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__clkbuf_1
X_4507_ BitStream_buffer.BS_buffer\[20\] _3048_ _3050_ BitStream_buffer.BS_buffer\[21\]
+ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__a22o_1
X_4438_ _2724_ _2800_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__nand2_1
X_4369_ _0761_ _2882_ _0638_ _2885_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__o22ai_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032__129 clknet_1_1__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6094__25 clknet_1_1__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__inv_2
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5995__95 clknet_1_0__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
X_3740_ BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__inv_2
XANTENNA_19 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3671_ _2831_ _2838_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
X_5410_ _1946_ _2117_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__or2_1
X_5341_ _2072_ _2055_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__and2_1
X_5272_ net7 BitStream_buffer.BS_buffer\[32\] _2024_ vssd1 vssd1 vccd1 vccd1 _2025_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4223_ _2751_ _2697_ _0431_ _2702_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__o22ai_1
X_4154_ _2856_ BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__nand2_1
X_4085_ _0516_ _3041_ _3043_ BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1
+ _0873_ sky130_fd_sc_hd__a22o_1
X_3105_ BitStream_buffer.BS_buffer\[74\] _2617_ BitStream_buffer.BS_buffer\[75\] _2624_
+ _2638_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4987_ _2870_ _2812_ _1763_ _1764_ _1765_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__o2111a_1
X_3938_ BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6070__3 clknet_1_1__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__inv_2
X_3869_ BitStream_buffer.BS_buffer\[22\] _0351_ BitStream_buffer.BS_buffer\[23\] _0354_
+ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__a221oi_1
X_5608_ net10 _2832_ _2229_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__mux2_1
X_5539_ _2208_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 exp_golomb_sel[0] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
XFILLER_0_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6015__113 clknet_1_0__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5890_ _2448_ _2507_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__nor2_1
X_4910_ BitStream_buffer.BS_buffer\[52\] _2948_ BitStream_buffer.BS_buffer\[53\] _2951_
+ _1689_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__a221oi_1
X_4841_ BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1 vccd1 _1622_
+ sky130_fd_sc_hd__inv_2
X_4772_ _0445_ _2807_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6061__155 clknet_1_0__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
X_3723_ BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3654_ BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3585_ _0363_ _0365_ _0366_ _0369_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5324_ _2060_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__clkbuf_4
X_5255_ _2011_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__inv_2
X_4206_ _0986_ _0988_ _0990_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5186_ _1959_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _2787_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ BitStream_buffer.BS_buffer\[44\] _2949_ BitStream_buffer.BS_buffer\[45\] _2952_
+ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5974__76 clknet_1_1__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__inv_2
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3370_ _2705_ _2774_ _2844_ _2903_ vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__and4_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _2910_ _0356_ _2914_ _0359_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__o22ai_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5942_ _2555_ _2557_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__nand2_1
X_5873_ _1310_ _2381_ _2490_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4824_ _0358_ _3061_ _0660_ _0322_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4755_ _0456_ _2734_ _2811_ _2738_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ BitStream_buffer.BS_buffer\[41\] _2949_ BitStream_buffer.BS_buffer\[42\] _2952_
+ _0496_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__a221oi_1
X_4686_ _2891_ BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3637_ BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3568_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5307_ _2048_ _2034_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__and2_1
X_6287_ net89 _0302_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[4\] sky130_fd_sc_hd__dfxtp_1
X_3499_ _3032_ _2672_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__nor2_2
X_5238_ _1997_ _1990_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__nand2_1
X_5169_ BitStream_buffer.buffer_index\[5\] vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2593_ clknet_0__2593_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2593_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4540_ _1313_ _1317_ _1320_ _1322_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__and4_1
X_4471_ _0638_ _2849_ _1252_ _1253_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3422_ BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__inv_2
X_6210_ net172 _0225_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[66\] sky130_fd_sc_hd__dfxtp_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3353_ BitStream_buffer.BS_buffer\[126\] _2876_ BitStream_buffer.BS_buffer\[127\]
+ _2879_ _2886_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__a221oi_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _2777_ _2672_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__nor2_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ BitStream_buffer.BS_buffer\[69\] _2991_ BitStream_buffer.BS_buffer\[70\] _2994_
+ _1801_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6067__161 clknet_1_1__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
X_5925_ _2522_ _2491_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5856_ _2421_ _2447_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4807_ _2640_ _2966_ _0508_ _2969_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5787_ _2402_ _2403_ _2408_ _2411_ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__o211ai_1
X_4738_ _0672_ _1517_ _1519_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4669_ _2814_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3971_ _0755_ _0757_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5710_ _2334_ _1310_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5641_ _2279_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5572_ _2231_ _2216_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4523_ _1275_ _1285_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__nor3_1
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4454_ _2898_ _2780_ _1235_ _1236_ _1237_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__o2111a_1
X_4385_ BitStream_buffer.BS_buffer\[47\] _2949_ BitStream_buffer.BS_buffer\[48\] _2952_
+ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__a221oi_1
X_3405_ BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__inv_2
X_3336_ BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__inv_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _1739_ _1754_ _1771_ _1784_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__and4_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _2799_ _2800_ vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__nand2_1
X_3198_ _2731_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5908_ _2489_ _2495_ _2522_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__nand3_1
X_5839_ BitStream_buffer.BitStream_buffer_output\[12\] _2432_ vssd1 vssd1 vccd1 vccd1
+ _2462_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4170_ BitStream_buffer.BS_buffer\[37\] _2929_ _2931_ BitStream_buffer.BS_buffer\[38\]
+ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__a22o_1
X_3121_ _2654_ _2621_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3954_ BitStream_buffer.BS_buffer\[35\] _2929_ _2931_ BitStream_buffer.BS_buffer\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3885_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__clkbuf_4
X_5624_ net7 BitStream_buffer.BS_buffer\[112\] _2267_ vssd1 vssd1 vccd1 vccd1 _2268_
+ sky130_fd_sc_hd__mux2_1
X_5555_ _2219_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5486_ _2170_ _2171_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__and2_1
X_4506_ _1286_ _1287_ _1288_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__or4_1
X_4437_ _2720_ _2804_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ BitStream_buffer.BS_buffer\[125\] _2863_ BitStream_buffer.BS_buffer\[126\]
+ _2866_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__a221oi_1
X_3319_ _2850_ _2852_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__or2_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _0646_ _3062_ _0523_ _0323_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__o22ai_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3670_ _0456_ _2813_ _0457_ _0458_ _0460_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__o2111a_1
X_5340_ net2 BitStream_buffer.BS_buffer\[21\] _2061_ vssd1 vssd1 vccd1 vccd1 _2072_
+ sky130_fd_sc_hd__mux2_1
X_5271_ _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4222_ _1006_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nor2_1
X_4153_ _0476_ _2852_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__or2_1
X_4084_ _0330_ _3034_ _3036_ _0325_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__a22o_1
X_3104_ _2625_ _2630_ _2631_ _2637_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4986_ _0481_ _2823_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__or2_1
X_3937_ _0476_ _2849_ _0723_ _0724_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3868_ _0657_ _0357_ _0534_ _0360_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__o22ai_1
X_3799_ _2819_ _2816_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__nand2_1
X_5607_ _2255_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
X_5538_ _2207_ _2195_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5469_ net6 BitStream_buffer.BS_buffer\[65\] _2157_ vssd1 vssd1 vccd1 vccd1 _2160_
+ sky130_fd_sc_hd__mux2_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 exp_golomb_sel[1] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _1577_ _1619_ _1620_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__nand3_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4771_ _2802_ _2838_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__nand2_1
X_3722_ _0512_ _3022_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3653_ _2788_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5323_ _2059_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3584_ _0370_ _0372_ _0373_ _0375_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5254_ net32 net31 vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__nand2_1
X_4205_ BitStream_buffer.BS_buffer\[33\] _0379_ BitStream_buffer.BS_buffer\[34\] _0383_
+ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__a221oi_1
X_5185_ _1958_ _1952_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__and2_1
X_4136_ _2888_ _2784_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__or2_1
X_4067_ _2939_ _2955_ _2942_ _2959_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4969_ _0694_ _2752_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6136__63 clknet_1_0__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__inv_2
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5941_ _2608_ _2556_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5872_ _2381_ BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1 vccd1
+ _2490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4823_ _0345_ _3054_ _0657_ _3057_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4754_ _0450_ _2712_ _1532_ _1533_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__o2111a_1
X_3705_ _0495_ _2955_ _2953_ _2959_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4685_ _0330_ _2875_ _0325_ _2879_ _1466_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__a221oi_1
X_3636_ _0423_ _2713_ _0424_ _0425_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3567_ _3028_ _0338_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__nand2_2
X_6286_ net88 _0301_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[5\] sky130_fd_sc_hd__dfxtp_1
X_5306_ net11 BitStream_buffer.BS_buffer\[43\] _2023_ vssd1 vssd1 vccd1 vccd1 _2048_
+ sky130_fd_sc_hd__mux2_1
X_5237_ _1995_ _2708_ _3012_ _1996_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__a31o_1
X_3498_ _3019_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5168_ BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__inv_2
X_5099_ _2855_ _0330_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__nand2_1
X_4119_ BitStream_buffer.BS_buffer\[83\] _2689_ _2766_ _2693_ _0905_ vssd1 vssd1 vccd1
+ vccd1 _0906_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6044__140 clknet_1_1__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2592_ clknet_0__2592_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2592_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _2859_ _0400_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__nand2_1
X_3421_ _2954_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__buf_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115__44 clknet_1_1__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__inv_2
X_3352_ _2880_ _2882_ _2883_ _2885_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__o22ai_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3283_ _2815_ _2816_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__nand2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6130__58 clknet_1_0__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__inv_2
X_5022_ _2631_ _2997_ _0556_ _3000_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__o22ai_1
X_5924_ _2328_ _2351_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__nand2_1
X_5855_ _2477_ _2417_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4806_ _1582_ _1584_ _1586_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__nand3b_1
X_5786_ _2348_ _2410_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4737_ _1518_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4668_ _2839_ _2796_ _1447_ _1448_ _1449_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__o2111a_1
X_3619_ _2650_ BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__nand2_1
X_4599_ BitStream_buffer.BS_buffer\[63\] _2981_ _2983_ BitStream_buffer.BS_buffer\[64\]
+ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__a22o_1
X_6269_ net71 _0284_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3970_ BitStream_buffer.BS_buffer\[63\] _3005_ BitStream_buffer.BS_buffer\[64\] _3008_
+ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _2278_ _2261_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5571_ net7 _2800_ _2230_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__mux2_1
X_4522_ _1296_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__nand2_1
X_4453_ _2791_ BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3404_ _2937_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__clkbuf_4
X_4384_ _2975_ _2955_ _0619_ _2959_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__o22ai_1
X_6123_ clknet_1_0__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__buf_1
X_3335_ _2868_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__buf_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__clkbuf_4
X_5005_ _1775_ _1777_ _1779_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__and4_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3197_ _2730_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__clkbuf_2
X_5907_ _2521_ _2523_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _2456_ _2460_ _2371_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__nand3_1
XFILLER_0_29_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5769_ BitStream_buffer.BitStream_buffer_output\[10\] BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3120_ _2653_ _2627_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__nor2_4
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3953_ BitStream_buffer.BS_buffer\[41\] _2924_ _2926_ BitStream_buffer.BS_buffer\[42\]
+ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3884_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5623_ _2266_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5554_ _2218_ _2216_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4505_ _0527_ _3041_ _3043_ _0650_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__a22o_1
X_5485_ _0404_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4436_ _2795_ _2717_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__or2_1
X_4367_ _2883_ _2869_ _2845_ _2872_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _2851_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__clkbuf_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _0660_ _3055_ _0537_ _3058_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__o22ai_1
X_3249_ _2620_ _2778_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5270_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ BitStream_buffer.BS_buffer\[76\] _2679_ _2682_ BitStream_buffer.BS_buffer\[77\]
+ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__a22o_1
X_4152_ _0926_ _0930_ _0934_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4083_ _3060_ _3026_ _3063_ _3030_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_37_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3103_ _2636_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__buf_6
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4985_ _2818_ BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3936_ _2859_ BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nand2_1
X_3867_ BitStream_buffer.BS_buffer\[25\] vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3798_ _2815_ _2792_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nand2_1
X_5606_ _2254_ _2240_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__and2_1
X_5537_ net16 _2762_ _2193_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__mux2_1
X_5468_ _2159_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
X_5399_ _2112_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
X_4419_ _0399_ BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__nand2_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 reset_n vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_4
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _2798_ _2781_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3721_ _3039_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3652_ _0427_ _0430_ _0436_ _0442_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__and4_1
X_3583_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5322_ BitStream_buffer.buffer_index\[6\] BitStream_buffer.buffer_index\[5\] _1947_
+ _1944_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__or4b_1
XFILLER_0_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5253_ _2009_ _2010_ _0675_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__a21oi_1
X_4204_ _2910_ _0386_ _2914_ _0390_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__o22ai_1
X_5184_ net4 _3044_ _1950_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__mux2_1
X_4135_ _0911_ _0913_ _0917_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4066_ BitStream_buffer.BS_buffer\[48\] _2935_ BitStream_buffer.BS_buffer\[49\] _2938_
+ _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4968_ _2748_ BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4899_ _2883_ _2889_ _1676_ _1677_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3919_ _2791_ _2781_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5940_ _2547_ _2371_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__nand2b_1
X_5871_ _2422_ _2488_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__nor2_1
X_4822_ BitStream_buffer.BS_buffer\[23\] _3047_ _3049_ BitStream_buffer.BS_buffer\[24\]
+ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4753_ _2723_ BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__nand2_1
X_3704_ BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4684_ _3024_ _2881_ _3027_ _2884_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3635_ _2724_ _2706_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__nand2_1
X_3566_ BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5305_ _2047_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
X_6285_ net87 _0300_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[6\] sky130_fd_sc_hd__dfxtp_1
X_3497_ _3024_ _3026_ _3027_ _3030_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__o22ai_1
X_5236_ BitStream_buffer.pc_previous\[6\] _2708_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5167_ _1938_ _1939_ net200 vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5098_ _3024_ _2851_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__or2_1
X_4118_ _0431_ _2697_ _2742_ _2702_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__o22ai_1
X_4049_ _2850_ _2869_ _0727_ _2872_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2591_ clknet_0__2591_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2591_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3420_ net36 _2907_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3351_ _2884_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__buf_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__clkbuf_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _1796_ _1797_ _1798_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5923_ _2537_ _2538_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5854_ _2473_ _2476_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__nand2_1
X_6028__125 clknet_1_0__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_0_63_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4805_ BitStream_buffer.BS_buffer\[51\] _2948_ BitStream_buffer.BS_buffer\[52\] _2951_
+ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__a221oi_1
X_5785_ _2321_ _2409_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__nand2_1
X_4736_ BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1 vccd1 _1518_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4667_ _2782_ _2807_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3618_ BitStream_buffer.BS_buffer\[75\] _2617_ BitStream_buffer.BS_buffer\[76\] _2624_
+ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__a221oi_1
X_4598_ _0505_ _2974_ _2996_ _2977_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__o22ai_1
X_3549_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6268_ net70 _0283_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dfxtp_1
X_5219_ _1981_ _1973_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__and2_1
X_6199_ net161 _0214_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[77\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5570_ _2229_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__clkbuf_4
X_4521_ _1298_ _1300_ _1302_ _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4452_ _2787_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__nand2_1
X_3403_ _2936_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4383_ BitStream_buffer.BS_buffer\[51\] _2935_ BitStream_buffer.BS_buffer\[52\] _2938_
+ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__a221oi_1
X_3334_ _2668_ _2847_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__nand2_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _2798_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__buf_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _2880_ _2889_ _1780_ _1781_ _1782_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__o2111a_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3196_ _2690_ _2711_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ _2522_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5837_ _2457_ _2459_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__nand2_1
X_5768_ _2361_ _2326_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__and2_1
X_4719_ _0660_ _3061_ _0537_ _0322_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5699_ _2312_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3952_ _0486_ _2916_ _2905_ _2920_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3883_ net19 vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5622_ _2265_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5553_ net11 _2714_ _2192_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4504_ _0770_ _3034_ _3036_ _3051_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5484_ net16 BitStream_buffer.BS_buffer\[70\] _2157_ vssd1 vssd1 vccd1 vccd1 _2170_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4435_ _1209_ _1213_ _1216_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4366_ _0512_ _2849_ _1148_ _1149_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__o2111a_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ net35 _2847_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__nand2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ BitStream_buffer.BS_buffer\[18\] _3048_ _3050_ BitStream_buffer.BS_buffer\[19\]
+ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__a22o_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _2781_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__inv_2
X_3179_ _2712_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__buf_2
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4220_ _0549_ _2670_ _0407_ _2675_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o22ai_1
X_4151_ _2870_ _2829_ _0935_ _0936_ _0937_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_49_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6085__17 clknet_1_0__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__inv_2
X_4082_ _0869_ _3022_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nor2_1
X_3102_ _2635_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4984_ _2814_ BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3935_ _2856_ BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__nand2_1
X_5986__87 clknet_1_1__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
XFILLER_0_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3866_ BitStream_buffer.BS_buffer\[26\] _0337_ BitStream_buffer.BS_buffer\[27\] _0341_
+ _0655_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__a221oi_1
X_5605_ net11 _2781_ _2229_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3797_ _2822_ _2797_ _0584_ _0585_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__o2111a_1
X_5536_ _2206_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5467_ _2158_ _2148_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__and2_1
X_4418_ _1171_ _1181_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__nor3_1
X_5398_ _0405_ BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__nand2_1
X_4349_ _2888_ _2780_ _1131_ _1132_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__o2111a_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3720_ _0504_ _0507_ _0510_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ _0437_ _2759_ _0438_ _0439_ _0441_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3582_ _2918_ _0338_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nand2_2
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5321_ _2058_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__clkbuf_1
X_5252_ _2001_ net28 vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__nand2_1
X_4203_ BitStream_buffer.BS_buffer\[21\] _0365_ BitStream_buffer.BS_buffer\[22\] _0369_
+ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a221oi_1
X_5183_ _1957_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4134_ _2737_ _2759_ _0918_ _0919_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__o2111a_1
X_4065_ _2972_ _2941_ _2975_ _2945_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _2745_ BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__nand2_1
X_4898_ _2880_ _2899_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__or2_1
X_3918_ _2787_ _2838_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3849_ _0638_ _3022_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__nor2_1
X_5519_ _0404_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5870_ _2459_ _2425_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4821_ _1598_ _1599_ _1600_ _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _2719_ BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4683_ _0400_ _2862_ BitStream_buffer.BS_buffer\[1\] _2866_ _1464_ vssd1 vssd1 vccd1
+ vccd1 _1465_ sky130_fd_sc_hd__a221oi_1
X_3703_ BitStream_buffer.BS_buffer\[45\] _2935_ BitStream_buffer.BS_buffer\[46\] _2938_
+ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3634_ _2720_ _2714_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3565_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__buf_2
X_6284_ net86 _0299_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[7\] sky130_fd_sc_hd__dfxtp_2
X_5304_ _2046_ _2034_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__and2_1
X_3496_ _3029_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__buf_4
X_5235_ _1994_ BitStream_buffer.pc_previous\[4\] BitStream_buffer.pc_previous\[5\]
+ BitStream_buffer.pc_previous\[6\] vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__a31o_1
X_5166_ _1941_ net199 vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2_1
X_5097_ _1862_ _1866_ _1870_ _1874_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__and4_1
X_4117_ _0902_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4048_ _0604_ _2849_ _0833_ _0834_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6005__104 clknet_1_0__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
XFILLER_0_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6051__146 clknet_1_0__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2590_ clknet_0__2590_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2590_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3350_ _2700_ _2847_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__nand2_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3281_ _2814_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__buf_2
X_5020_ BitStream_buffer.BS_buffer\[61\] _2985_ _2987_ BitStream_buffer.BS_buffer\[62\]
+ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__a22o_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5922_ _2447_ _2416_ _2475_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__nor3_1
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5853_ _2451_ _2448_ _2475_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5784_ BitStream_buffer.BitStream_buffer_output\[6\] BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__nand2_1
X_4804_ _0499_ _2954_ _2963_ _2958_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4735_ _1473_ _1515_ _1516_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__nand3_1
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ _2802_ _2832_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4597_ _3009_ _2967_ _0632_ _2970_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__o22ai_1
X_3617_ _0407_ _2630_ _2625_ _2637_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__o22ai_1
X_3548_ _0339_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__clkbuf_2
X_6267_ net69 _0282_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[32\] sky130_fd_sc_hd__dfxtp_2
X_3479_ _3012_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__inv_2
X_5218_ net8 _0521_ _1949_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__mux2_1
X_6198_ net160 _0213_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[78\] sky130_fd_sc_hd__dfxtp_2
X_5149_ _0622_ _0385_ _0495_ _0389_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_81_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4520_ BitStream_buffer.BS_buffer\[36\] _0379_ BitStream_buffer.BS_buffer\[37\] _0383_
+ _1303_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4451_ _2894_ _2784_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__or2_1
X_3402_ _2695_ _2907_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _0499_ _2941_ _2963_ _2945_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__o22ai_1
X_3333_ BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__inv_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _2777_ _2643_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__nor2_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5003_ _0476_ _2899_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__or2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _2728_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__buf_2
X_5905_ _2381_ _1414_ _1206_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__a21oi_2
X_6073__6 clknet_1_1__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__inv_2
XFILLER_0_48_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5836_ BitStream_buffer.BitStream_buffer_output\[6\] _2381_ _2458_ vssd1 vssd1 vccd1
+ vccd1 _2459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5767_ _2384_ _2391_ _2371_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__nand3_1
X_5698_ _2322_ _1622_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__nand2_1
X_4718_ _0657_ _3054_ _0534_ _3057_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4649_ _2795_ _2712_ _1428_ _1429_ _1430_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _0739_ _2909_ _0613_ _2912_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3882_ _2598_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__buf_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5621_ _1945_ _2118_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5552_ _2217_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4503_ _3053_ _3026_ _3056_ _3030_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5483_ _2169_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__clkbuf_1
X_4434_ _2762_ _2689_ _2756_ _2693_ _1217_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4365_ _2859_ BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__inv_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _1078_ _1079_ _1080_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__or4_1
X_6035_ clknet_1_1__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__buf_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__clkbuf_4
X_3178_ net35 _2711_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__nand2_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5819_ _2440_ _2441_ _2442_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4150_ _0481_ _2841_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or2_1
X_3101_ _2603_ _2634_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__or2_1
X_4081_ BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4983_ _2888_ _2796_ _1759_ _1760_ _1761_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3934_ _2883_ _2852_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3865_ _0654_ _0344_ _0531_ _0347_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5604_ _2253_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3796_ _2795_ _2808_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__or2_1
X_5535_ _2205_ _2195_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5466_ net7 BitStream_buffer.BS_buffer\[64\] _2157_ vssd1 vssd1 vccd1 vccd1 _2158_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ _1192_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__nand2_1
X_5397_ _2111_ _2101_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc\[3\] sky130_fd_sc_hd__xor2_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4348_ _2791_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nand2_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4279_ _0619_ _2955_ _0492_ _2959_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3650_ _0440_ _2771_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or2_1
X_3581_ BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5320_ _2057_ _2055_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__and2_1
X_5251_ _1998_ _1993_ _2008_ _2001_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4202_ _0534_ _0372_ _0355_ _0375_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__o22ai_1
X_5182_ _1956_ _1952_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__and2_1
X_4133_ _0423_ _2771_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _0848_ _0849_ _0850_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4966_ _2781_ _2728_ _2832_ _2731_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4897_ _0604_ _2895_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__or2_1
X_3917_ _0464_ _2784_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3848_ BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__inv_2
X_3779_ _0568_ _2735_ _0428_ _2739_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__o22ai_1
X_5518_ net7 BitStream_buffer.BS_buffer\[80\] _2193_ vssd1 vssd1 vccd1 vccd1 _2194_
+ sky130_fd_sc_hd__mux2_1
X_5449_ _2145_ _2127_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6127__55 clknet_1_1__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__inv_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142__69 clknet_1_1__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__inv_2
XFILLER_0_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4820_ _3051_ _3040_ _3042_ _0521_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4751_ _0459_ _2716_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4682_ _0604_ _2868_ _0476_ _2871_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__o22ai_1
X_3702_ _0492_ _2941_ _2939_ _2945_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3633_ _2737_ _2717_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3564_ _2680_ _0338_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__nand2_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5303_ net12 BitStream_buffer.BS_buffer\[42\] _2023_ vssd1 vssd1 vccd1 vccd1 _2046_
+ sky130_fd_sc_hd__mux2_1
X_6283_ net85 _0298_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[8\] sky130_fd_sc_hd__dfxtp_1
X_3495_ _3028_ _3020_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__nand2_2
X_5234_ BitStream_buffer.pc_previous\[1\] BitStream_buffer.pc_previous\[0\] BitStream_buffer.pc_previous\[2\]
+ BitStream_buffer.pc_previous\[3\] vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__and4_1
X_5165_ net198 net29 vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4116_ BitStream_buffer.BS_buffer\[75\] _2679_ _2682_ BitStream_buffer.BS_buffer\[76\]
+ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__a22o_1
X_5096_ _2880_ _2828_ _1871_ _1872_ _1873_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__o2111a_1
X_4047_ _2859_ BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4949_ _0440_ _2629_ _2769_ _2636_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970__72 clknet_1_1__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__inv_2
XFILLER_0_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _2777_ _2677_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__nor2_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5921_ _2536_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5852_ _2474_ _2415_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5783_ _2352_ _2353_ _2407_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__nand3_1
X_4803_ BitStream_buffer.BS_buffer\[55\] _2934_ BitStream_buffer.BS_buffer\[56\] _2937_
+ _1583_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__a221oi_1
X_4734_ _0398_ _0527_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4665_ _2798_ _2788_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4596_ _1374_ _1376_ _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__nand3b_1
X_3616_ BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
X_6106__36 clknet_1_1__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__inv_2
X_3547_ _2628_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__and2_1
X_6266_ net68 _0281_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[33\] sky130_fd_sc_hd__dfxtp_4
X_3478_ _2690_ _2965_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__nand2_2
X_5217_ _1980_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__clkbuf_1
X_6197_ net159 _0212_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[79\] sky130_fd_sc_hd__dfxtp_2
X_5148_ _0387_ _0364_ BitStream_buffer.BS_buffer\[31\] _0368_ _1925_ vssd1 vssd1 vccd1
+ vccd1 _1926_ sky130_fd_sc_hd__a221oi_1
X_5079_ _2822_ _2758_ _1854_ _1855_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4450_ _1223_ _1225_ _1229_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4381_ _1162_ _1163_ _1164_ _1165_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__or4_1
X_3401_ _2934_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3332_ _2865_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__buf_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _2796_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__buf_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034__131 clknet_1_1__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
X_5002_ _0730_ _2895_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__or2_1
X_3194_ _2710_ _2687_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__nor2_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5904_ _2493_ _2453_ _2495_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5835_ _2368_ _1622_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__nand2_1
X_5766_ _2387_ _2390_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5697_ BitStream_buffer.BitStream_buffer_output\[7\] _2321_ vssd1 vssd1 vccd1 vccd1
+ _2322_ sky130_fd_sc_hd__nor2_1
X_4717_ BitStream_buffer.BS_buffer\[22\] _3047_ _3049_ BitStream_buffer.BS_buffer\[23\]
+ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4648_ _2723_ _2804_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4579_ _3027_ _2882_ _0869_ _2885_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__o22ai_1
X_6249_ net51 _0264_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[18\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3950_ BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__inv_2
X_3881_ BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1 vccd1 vccd1 _0671_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5620_ _2264_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
X_5551_ _2215_ _2216_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__and2_1
X_4502_ _0640_ _3022_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5482_ _2168_ _2148_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4433_ _2769_ _2697_ _0434_ _2702_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__o22ai_1
X_4364_ _2856_ BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__nand2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _2848_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__clkbuf_4
X_4295_ _0330_ _3041_ _3043_ _0325_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__a22o_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _2779_ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__clkbuf_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3177_ _2710_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5818_ _2354_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5749_ _2373_ _2607_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3100_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4080_ _0863_ _0865_ _0867_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__nand3b_1
X_4982_ _0464_ _2807_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3933_ _0709_ _0713_ _0717_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__and4_1
X_3864_ _0380_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5603_ _2252_ _2240_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3795_ _2803_ _2820_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__nand2_1
X_5534_ net2 _2768_ _2193_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5465_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4416_ _1194_ _1196_ _1198_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__and4_1
X_5396_ _2110_ _2103_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__and2b_2
X_4347_ _2787_ BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__nand2_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4278_ BitStream_buffer.BS_buffer\[50\] _2935_ BitStream_buffer.BS_buffer\[51\] _2938_
+ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a221oi_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _2761_ _2762_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3580_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5250_ net28 _1943_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__or2_1
X_4201_ BitStream_buffer.BS_buffer\[25\] _0351_ BitStream_buffer.BS_buffer\[26\] _0354_
+ _0987_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__a221oi_1
X_5181_ net5 _3039_ _1950_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__mux2_1
X_4132_ _2765_ _2706_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4063_ BitStream_buffer.BS_buffer\[36\] _2929_ _2931_ BitStream_buffer.BS_buffer\[37\]
+ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4965_ _0444_ _2734_ _2775_ _2738_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__o22ai_1
X_3916_ _0693_ _0696_ _0700_ _0704_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4896_ _2891_ BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3847_ _0631_ _0634_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__inv_2
X_5517_ _2192_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5448_ net11 BitStream_buffer.BS_buffer\[59\] _2120_ vssd1 vssd1 vccd1 vccd1 _2145_
+ sky130_fd_sc_hd__mux2_1
X_5379_ BitStream_buffer.pc_previous\[2\] BitStream_buffer.exp_golomb_len\[2\] vssd1
+ vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2589_ clknet_0__2589_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2589_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750_ _1521_ _1525_ _1528_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4681_ _0869_ _2848_ _1460_ _1461_ _1462_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__o2111a_1
X_3701_ BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3632_ _2721_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3563_ BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__inv_2
X_5302_ _2045_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6282_ net84 _0297_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[9\] sky130_fd_sc_hd__dfxtp_1
X_3494_ _2677_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__inv_2
X_5233_ BitStream_buffer.pc\[6\] _1948_ _1990_ _1992_ vssd1 vssd1 vccd1 vccd1 _1993_
+ sky130_fd_sc_hd__a31oi_2
X_5164_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__inv_2
X_4115_ _0407_ _2670_ _2625_ _2675_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__o22ai_1
X_5095_ _2845_ _2840_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__or2_1
X_4046_ _2856_ BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4948_ _0672_ _1725_ _1727_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__o21a_1
X_4879_ _2814_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5920_ _2529_ _2415_ _2503_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5851_ _2461_ _2471_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__nand2_1
X_5782_ _2405_ _2406_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4802_ _2999_ _2940_ _0858_ _2944_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4733_ _1483_ _1493_ _1514_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__nor3_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4664_ _2894_ _2779_ _1443_ _1444_ _1445_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__o2111a_1
X_3615_ _2599_ _0402_ _0406_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4595_ BitStream_buffer.BS_buffer\[49\] _2949_ BitStream_buffer.BS_buffer\[50\] _2952_
+ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__a221oi_1
X_3546_ _0334_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__clkbuf_4
X_6265_ net67 _0280_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[34\] sky130_fd_sc_hd__dfxtp_2
X_5216_ _1979_ _1973_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__and2_1
X_3477_ _3010_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6196_ net158 _0211_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[80\] sky130_fd_sc_hd__dfxtp_2
X_5147_ _0663_ _0371_ _0540_ _0374_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__o22ai_1
X_5078_ _2795_ _2770_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__or2_1
X_6011__110 clknet_1_1__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
X_4029_ _2787_ _2836_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4380_ BitStream_buffer.BS_buffer\[39\] _2929_ _2931_ BitStream_buffer.BS_buffer\[40\]
+ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__a22o_1
X_3400_ _2922_ _2699_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__nor2_2
X_3331_ _2864_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__clkbuf_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _2659_ _2778_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__nand2_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _2891_ BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__nand2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _2707_ _2713_ _2718_ _2722_ _2726_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5903_ _2518_ _2519_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5834_ _2370_ _2390_ _2425_ vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5765_ _2388_ _2389_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5696_ _2320_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__inv_2
X_4716_ _1494_ _1495_ _1496_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4647_ _2719_ _2820_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__nand2_1
X_4578_ _0400_ _2865_ BitStream_buffer.BS_buffer\[127\] _2863_ _1360_ vssd1 vssd1
+ vccd1 vccd1 _1361_ sky130_fd_sc_hd__a221oi_1
X_3529_ BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__inv_2
X_6248_ net50 _0263_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[19\] sky130_fd_sc_hd__dfxtp_2
X_6179_ net141 _0194_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[97\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018__116 clknet_1_1__leaf__2586_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
X_6097__28 clknet_1_0__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__inv_2
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998__98 clknet_1_1__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6064__158 clknet_1_0__leaf__2590_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
X_3880_ _0612_ _0668_ _0669_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5550_ net19 vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__clkbuf_2
X_5481_ net2 BitStream_buffer.BS_buffer\[69\] _2157_ vssd1 vssd1 vccd1 vccd1 _2168_
+ sky130_fd_sc_hd__mux2_1
X_4501_ _1280_ _1282_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4432_ _1214_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4363_ _0730_ _2852_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__or2_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _0527_ _3034_ _3036_ _0650_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__a22o_1
X_3314_ _2620_ _2847_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__nand2_2
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ net35 _2778_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__nand2_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _2709_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5817_ BitStream_buffer.BitStream_buffer_output\[9\] _2405_ vssd1 vssd1 vccd1 vccd1
+ _2441_ sky130_fd_sc_hd__nor2_1
X_5748_ _2359_ _2365_ _2372_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__nand3_2
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ _2304_ _2285_ _2117_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4981_ _2802_ BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__nand2_1
X_3932_ _0481_ _2829_ _0718_ _0719_ _0720_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3863_ _0644_ _0652_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__nor2_1
X_5602_ net12 _2788_ _2229_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__mux2_1
X_3794_ _2799_ _2804_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__nand2_1
X_5533_ _2204_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _1944_ _1991_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__nand2_4
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5395_ BitStream_buffer.pc_previous\[3\] BitStream_buffer.exp_golomb_len\[3\] vssd1
+ vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__nor2_1
X_4415_ BitStream_buffer.BS_buffer\[35\] _0379_ BitStream_buffer.BS_buffer\[36\] _0383_
+ _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__a221oi_1
X_4346_ _0481_ _2784_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__or2_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4277_ _2963_ _2941_ _2968_ _2945_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__o22ai_1
X_3228_ BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__clkbuf_4
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ _2692_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5977__79 clknet_1_0__leaf__2582_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__inv_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6047__142 clknet_1_0__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4200_ _0531_ _0357_ _0342_ _0360_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__o22ai_1
X_5180_ _1955_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__clkbuf_1
X_4131_ _2761_ _2714_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__nand2_1
X_4062_ BitStream_buffer.BS_buffer\[42\] _2924_ _2926_ BitStream_buffer.BS_buffer\[43\]
+ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4964_ _0459_ _2712_ _1740_ _1741_ _1742_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3915_ _0423_ _2759_ _0701_ _0702_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4895_ _0527_ _2875_ _0650_ _2878_ _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3846_ BitStream_buffer.BS_buffer\[62\] _3005_ BitStream_buffer.BS_buffer\[63\] _3008_
+ _0635_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3777_ _2715_ _2713_ _0564_ _0565_ _0566_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__o2111a_1
X_5516_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__buf_2
X_5447_ _2144_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
X_5378_ BitStream_buffer.pc_previous\[2\] BitStream_buffer.exp_golomb_len\[2\] vssd1
+ vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__or2_1
X_4329_ _2768_ _2689_ _2762_ _2693_ _1113_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2588_ clknet_0__2588_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2588_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3700_ _0487_ _0488_ _0489_ _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4680_ _2858_ _3039_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3631_ _0409_ _0414_ _0418_ _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and4_1
X_3562_ _0353_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__clkbuf_4
X_5301_ _2044_ _2034_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__and2_1
X_6281_ net83 _0296_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[10\] sky130_fd_sc_hd__dfxtp_1
X_3493_ BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5232_ _3012_ _2708_ _1990_ _1991_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__and4_1
X_5163_ net30 net29 vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__nor2_1
X_4114_ _2664_ _2646_ _0898_ _0899_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__o2111a_1
X_5094_ _2834_ BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__nand2_1
X_4045_ _2880_ _2852_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4947_ _1726_ _2598_ _0674_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4878_ _2827_ _2796_ _1655_ _1656_ _1657_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3829_ BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6132__60 clknet_1_0__leaf__2596_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__inv_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5850_ _2452_ _2472_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5781_ BitStream_buffer.BitStream_buffer_output\[8\] BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__nand2_1
X_4801_ _1578_ _1579_ _1580_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__or4_1
X_4732_ _1504_ _1513_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4663_ _2790_ BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__nand2_1
X_3614_ BitStream_buffer.BitStream_buffer_output\[15\] _0403_ _0405_ vssd1 vssd1 vccd1
+ vccd1 _0406_ sky130_fd_sc_hd__o21a_1
X_4594_ _2968_ _2955_ _2972_ _2959_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__o22ai_1
X_3545_ _0336_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__buf_2
X_6264_ net66 _0279_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[35\] sky130_fd_sc_hd__dfxtp_2
X_3476_ _2943_ _2965_ vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5215_ net9 _3051_ _1949_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6195_ net157 _0210_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[81\] sky130_fd_sc_hd__dfxtp_2
X_5146_ BitStream_buffer.BS_buffer\[34\] _0350_ BitStream_buffer.BS_buffer\[35\] _0353_
+ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__a221oi_1
X_5077_ _2764_ _2804_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__nand2_1
X_4028_ _2827_ _2784_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3330_ _2680_ _2847_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__and2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _0650_ _2875_ _0770_ _2878_ _1778_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__a221oi_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__inv_2
X_6111__41 clknet_1_0__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__inv_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _2724_ _2725_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5902_ _2504_ _2511_ _2375_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__o21ai_1
X_5833_ _2453_ _2425_ _2455_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__nand3_1
XFILLER_0_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5764_ _2361_ _1830_ _2328_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6041__137 clknet_1_1__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
X_5695_ BitStream_buffer.BitStream_buffer_output\[6\] BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__nor2_1
X_4715_ _0770_ _3040_ _3042_ _3051_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4646_ _2822_ _2716_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4577_ _0476_ _2869_ _2880_ _2872_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3528_ _3061_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__buf_2
X_6247_ net49 _0262_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[20\] sky130_fd_sc_hd__dfxtp_2
X_3459_ _2628_ _2965_ vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__and2_1
X_6178_ net140 _0193_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[98\] sky130_fd_sc_hd__dfxtp_1
X_5129_ _2698_ _3010_ BitStream_buffer.BS_buffer\[77\] _3013_ vssd1 vssd1 vccd1 vccd1
+ _1907_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5480_ _2167_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4500_ BitStream_buffer.BS_buffer\[68\] _3005_ BitStream_buffer.BS_buffer\[69\] _3008_
+ _1283_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _1171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4431_ BitStream_buffer.BS_buffer\[78\] _2679_ _2682_ BitStream_buffer.BS_buffer\[79\]
+ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__a22o_1
X_4362_ _1134_ _1138_ _1142_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__and4_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ clknet_1_1__leaf__2580_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__buf_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _0648_ _3026_ _0525_ _3030_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__o22ai_1
X_3313_ _2846_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__clkbuf_4
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _2777_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__inv_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ BitStream_buffer.pc\[5\] _2708_ _2600_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__or3_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5816_ _1102_ _2404_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5747_ _2370_ _2371_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5678_ BitStream_buffer.buffer_index\[4\] _1944_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__or2_1
X_4629_ _0399_ _0325_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4980_ _2798_ _2838_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__nand2_1
X_3931_ _2888_ _2841_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__or2_1
X_3862_ _0645_ _0647_ _0649_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__or4_1
X_5601_ _2251_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
X_5532_ _2203_ _2195_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__and2_1
X_3793_ _2782_ _2780_ _0580_ _0581_ _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5463_ _2155_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5394_ _2109_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__inv_2
X_4414_ _0486_ _0386_ _2905_ _0390_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4345_ _1119_ _1121_ _1125_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__and4_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4276_ _1058_ _1059_ _1060_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__or4_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _2760_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__buf_2
X_3158_ _2691_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__clkbuf_2
X_3089_ _2622_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6139__66 clknet_1_1__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__inv_2
XFILLER_0_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4130_ _0440_ _2744_ _0914_ _0915_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__o2111a_1
X_4061_ _0613_ _2916_ _0486_ _2920_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6081__13 clknet_1_0__leaf__2592_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__inv_2
X_4963_ _2723_ BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3914_ _0437_ _2771_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__or2_1
X_4894_ _0640_ _2881_ _0514_ _2884_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_61_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5982__83 clknet_1_1__leaf__2583_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__inv_2
X_3845_ _2640_ _3011_ BitStream_buffer.BS_buffer\[65\] _3014_ vssd1 vssd1 vccd1 vccd1
+ _0635_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3776_ _2724_ _2721_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__nand2_1
X_5515_ _1945_ BitStream_buffer.buffer_index\[5\] _1947_ _1944_ vssd1 vssd1 vccd1
+ vccd1 _2191_ sky130_fd_sc_hd__or4b_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ _2143_ _2127_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__and2_1
X_5377_ _2611_ _2097_ _2096_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__o21ai_4
X_4328_ _0434_ _2697_ _2751_ _2702_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__o22ai_1
X_4259_ _2856_ _0400_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2587_ clknet_0__2587_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2587_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ BitStream_buffer.BS_buffer\[79\] _2689_ BitStream_buffer.BS_buffer\[80\] _2693_
+ _0420_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__a221oi_1
X_3561_ _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__clkbuf_2
X_5300_ net13 BitStream_buffer.BS_buffer\[41\] _2024_ vssd1 vssd1 vccd1 vccd1 _2044_
+ sky130_fd_sc_hd__mux2_1
X_6118__47 clknet_1_0__leaf__2595_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__inv_2
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6280_ net82 _0295_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[11\] sky130_fd_sc_hd__dfxtp_1
X_3492_ _3025_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__buf_4
X_5231_ _1946_ _1947_ BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 _1991_
+ sky130_fd_sc_hd__and3_1
X_5162_ _1937_ _1936_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__and2_1
X_5093_ _2830_ BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__nand2_1
X_4113_ _2631_ _2661_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__or2_1
X_6076__9 clknet_1_0__leaf__2591_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__inv_2
X_4044_ _0819_ _0823_ _0827_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4946_ BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1 vccd1 _1726_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4877_ _2839_ _2807_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__or2_1
X_3828_ _0614_ _0615_ _0616_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3759_ BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__inv_2
X_5429_ _2132_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4800_ BitStream_buffer.BS_buffer\[43\] _2928_ _2930_ BitStream_buffer.BS_buffer\[44\]
+ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__a22o_1
X_5780_ _2404_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4731_ _1506_ _1508_ _1510_ _1512_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4662_ _2786_ BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3613_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4593_ BitStream_buffer.BS_buffer\[53\] _2935_ BitStream_buffer.BS_buffer\[54\] _2938_
+ _1375_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__a221oi_1
X_3544_ _0335_ _2634_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nor2_2
XFILLER_0_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6263_ net65 _0278_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[36\] sky130_fd_sc_hd__dfxtp_2
X_3475_ BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5214_ _1978_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6194_ net156 _0209_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[82\] sky130_fd_sc_hd__dfxtp_2
X_5145_ _2905_ _0356_ _2910_ _0359_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5076_ _2760_ _2820_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__nand2_1
X_4027_ _0804_ _0806_ _0810_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4929_ _0355_ _3061_ _0358_ _0322_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2589_ _2589_ vssd1 vssd1 vccd1 vccd1 clknet_0__2589_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _2775_ _2780_ _2785_ _2789_ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__o2111a_1
X_3191_ BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__buf_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5901_ _2508_ _2374_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5832_ _1414_ _2381_ _2454_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5763_ _2329_ _2360_ _1622_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4714_ _0521_ _3033_ _3035_ BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1
+ _1496_ sky130_fd_sc_hd__a22o_1
X_5694_ _2312_ _2318_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4645_ _1417_ _1421_ _1424_ _1426_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4576_ _0761_ _2849_ _1356_ _1357_ _1358_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__o2111a_1
X_3527_ net36 _3020_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__nand2_2
X_6246_ net48 _0261_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[21\] sky130_fd_sc_hd__dfxtp_2
X_3458_ _2991_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__clkbuf_4
X_3389_ _2922_ _2677_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__nor2_2
X_6177_ net139 _0192_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[99\] sky130_fd_sc_hd__dfxtp_2
X_5128_ BitStream_buffer.BS_buffer\[70\] _2991_ BitStream_buffer.BS_buffer\[71\] _2994_
+ _1905_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__a221oi_1
X_5059_ _0419_ _2645_ _1834_ _1835_ _1836_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4430_ _2694_ _2670_ _2698_ _2675_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__o22ai_1
XANTENNA_2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4361_ _0473_ _2829_ _1143_ _1144_ _1145_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _3024_ _3022_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nor2_1
X_3312_ BitStream_buffer.pc\[6\] BitStream_buffer.pc\[4\] BitStream_buffer.pc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__and3_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _2776_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__clkbuf_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5815_ _2314_ _2438_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5746_ _2345_ _2329_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__nor2_2
X_5677_ _2303_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4628_ _1379_ _1389_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nor3_1
X_4559_ _0481_ _2780_ _1339_ _1340_ _1341_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__o2111a_1
X_6229_ net191 _0244_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc_previous\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _2835_ BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3861_ _0650_ _0327_ _0329_ _0527_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3792_ _2791_ _2788_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__nand2_1
X_5600_ _2250_ _2240_ vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__and2_1
X_5531_ net3 _2766_ _2193_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5462_ _2154_ _2148_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5393_ _0405_ BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__nand2_1
X_4413_ BitStream_buffer.BS_buffer\[23\] _0365_ BitStream_buffer.BS_buffer\[24\] _0369_
+ _1197_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__a221oi_1
X_4344_ _0428_ _2759_ _1126_ _1127_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__o2111a_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4275_ BitStream_buffer.BS_buffer\[38\] _2929_ _2931_ BitStream_buffer.BS_buffer\[39\]
+ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__a22o_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _2710_ _2677_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__nor2_2
X_3157_ _2690_ _2602_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3088_ _2620_ _2621_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5729_ _2352_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4060_ _0847_ _2909_ _0739_ _2912_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__o22ai_1
X_4962_ _2719_ BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4893_ _3039_ _2862_ _3044_ _2865_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__a221oi_1
X_3913_ _2765_ _2756_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3844_ BitStream_buffer.BS_buffer\[58\] _2992_ BitStream_buffer.BS_buffer\[59\] _2995_
+ _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3775_ _2720_ _2736_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5514_ _2190_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
X_5445_ net12 BitStream_buffer.BS_buffer\[58\] _2120_ vssd1 vssd1 vccd1 vccd1 _2143_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5376_ _2095_ _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__nand2_2
X_4327_ _1110_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nor2_1
X_4258_ _0604_ _2852_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__or2_1
X_3209_ _2654_ _2711_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__nand2_2
X_4189_ _0325_ _3034_ _3036_ _0527_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2586_ clknet_0__2586_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2586_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3560_ _2668_ _0338_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5230_ net28 _1941_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__nor2_1
X_3491_ _2680_ _3020_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__nand2_2
X_5161_ _1936_ _1937_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5092_ _2867_ _2812_ _1867_ _1868_ _1869_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__o2111a_1
X_4112_ _0415_ _2656_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__or2_1
X_4043_ _2894_ _2829_ _0828_ _0829_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4945_ _1681_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4876_ _2802_ _2836_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__nand2_1
X_3827_ BitStream_buffer.BS_buffer\[34\] _2929_ _2931_ BitStream_buffer.BS_buffer\[35\]
+ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3758_ _2599_ _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__o21a_1
X_3689_ _2870_ _2896_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__or2_1
X_5428_ _2131_ _2127_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__and2_1
X_5359_ net11 BitStream_buffer.BS_buffer\[27\] _2060_ vssd1 vssd1 vccd1 vccd1 _2085_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4730_ BitStream_buffer.BS_buffer\[38\] _0378_ BitStream_buffer.BS_buffer\[39\] _0383_
+ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4661_ _2867_ _2783_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3612_ net19 vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4592_ _0750_ _2941_ _0626_ _2945_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__o22ai_1
X_3543_ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
X_6262_ net64 _0277_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[37\] sky130_fd_sc_hd__dfxtp_2
X_3474_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__clkbuf_4
X_6193_ net155 _0208_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[83\] sky130_fd_sc_hd__dfxtp_2
X_5213_ _1977_ _1973_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__and2_1
X_5144_ BitStream_buffer.BS_buffer\[38\] _0336_ BitStream_buffer.BS_buffer\[39\] _0340_
+ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__a221oi_1
X_5075_ _0568_ _2743_ _1850_ _1851_ _1852_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4026_ _2715_ _2759_ _0811_ _0812_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4928_ _0342_ _3054_ _0345_ _3057_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4859_ _2822_ _2712_ _1636_ _1637_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__o2111a_1
Xclkbuf_0__2588_ _2588_ vssd1 vssd1 vccd1 vccd1 clknet_0__2588_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _2723_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__buf_4
X_5900_ _2509_ _2515_ _2517_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__o21ai_2
X_5831_ _2381_ BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1 vccd1
+ _2454_ sky130_fd_sc_hd__nand2_1
X_5762_ _2385_ _2386_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4713_ _0646_ _3025_ _0523_ _3029_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__o22ai_1
X_5693_ _2317_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__inv_2
X_4644_ _2725_ _2688_ _2706_ _2692_ _1425_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4575_ _2859_ BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nand2_1
X_3526_ BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__inv_2
X_6245_ net47 _0260_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[22\] sky130_fd_sc_hd__dfxtp_2
X_3457_ _2979_ _2634_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__nor2_2
X_6102__32 clknet_1_1__leaf__2594_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__inv_2
X_3388_ _2906_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__inv_2
X_6176_ net138 _0191_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[100\] sky130_fd_sc_hd__dfxtp_1
X_5127_ _2625_ _2997_ _2631_ _3000_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__o22ai_1
X_5058_ _2742_ _2660_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__or2_1
X_4009_ _0795_ _0796_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6001__101 clknet_1_1__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
XANTENNA_3 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4360_ _2870_ _2841_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__or2_1
X_3311_ BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__inv_2
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _1072_ _1074_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nand3b_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ BitStream_buffer.pc\[4\] _2708_ _2601_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__or3_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _2706_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5814_ _2313_ BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1 vccd1 vccd1
+ _2438_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5745_ _2367_ _2369_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5676_ _2118_ _2285_ _2302_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__and3_1
X_4627_ _1400_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4558_ _2791_ BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__nand2_1
X_3509_ _3042_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__clkbuf_4
X_4489_ _2972_ _2955_ _2975_ _2959_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__o22ai_1
X_6228_ net190 _0243_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[48\] sky130_fd_sc_hd__dfxtp_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ net121 _0174_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[117\] sky130_fd_sc_hd__dfxtp_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3860_ BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3791_ _2787_ _2832_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__nand2_1
X_5530_ _2202_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5461_ net1 BitStream_buffer.BS_buffer\[63\] _2120_ vssd1 vssd1 vccd1 vccd1 _2154_
+ sky130_fd_sc_hd__mux2_1
X_4412_ _0345_ _0372_ _0657_ _0375_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__o22ai_1
X_5392_ BitStream_buffer.pc_previous\[4\] _2104_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.pc\[4\]
+ sky130_fd_sc_hd__xor2_4
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4343_ _2737_ _2771_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4274_ BitStream_buffer.BS_buffer\[44\] _2924_ _2926_ BitStream_buffer.BS_buffer\[45\]
+ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__a22o_1
X_6013_ clknet_1_1__leaf__2581_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__buf_1
X_3225_ _2758_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__buf_2
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3156_ _2685_ _2619_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__nor2_4
X_3087_ _2602_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6008__107 clknet_1_0__leaf__2585_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5728_ _2341_ _2346_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__nand2_2
X_3989_ _0358_ _0372_ _0660_ _0375_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5659_ _2291_ _2285_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6054__149 clknet_1_1__leaf__2589_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6145__1 clknet_1_1__leaf__2581_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__inv_2
X_4961_ _0456_ _2716_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__or2_1
X_3912_ _2761_ _2706_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__nand2_1
X_4892_ _3018_ _2868_ _0730_ _2871_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3843_ _0632_ _2998_ _0505_ _3001_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__o22ai_1
X_3774_ _2733_ _2717_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5513_ _2189_ _2171_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__and2_1
X_5444_ _2142_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6144__71 clknet_1_1__leaf__2597_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__inv_2
XFILLER_0_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5375_ BitStream_buffer.pc_previous\[1\] BitStream_buffer.exp_golomb_len\[1\] vssd1
+ vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__nand2_1
X_4326_ BitStream_buffer.BS_buffer\[77\] _2679_ _2682_ BitStream_buffer.BS_buffer\[78\]
+ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__a22o_1
X_4257_ _1030_ _1034_ _1038_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__and4_1
X_4188_ _0525_ _3026_ _3060_ _3030_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__o22ai_1
X_3208_ BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__inv_2
X_3139_ _2672_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2585_ clknet_0__2585_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2585_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3490_ BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6037__133 clknet_1_0__leaf__2588_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
X_5160_ net33 net32 vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__nor2_1
X_5091_ _2894_ _2823_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__or2_1
X_4111_ _2650_ BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__nand2_1
X_4042_ _2898_ _2841_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4944_ _0398_ _0770_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4875_ _2798_ _2832_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3826_ BitStream_buffer.BS_buffer\[40\] _2924_ _2926_ BitStream_buffer.BS_buffer\[41\]
+ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3757_ BitStream_buffer.BitStream_buffer_output\[14\] _0403_ _0405_ vssd1 vssd1 vccd1
+ vccd1 _0548_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3688_ _2892_ BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__nand2_1
X_5427_ net3 BitStream_buffer.BS_buffer\[52\] _2121_ vssd1 vssd1 vccd1 vccd1 _2131_
+ sky130_fd_sc_hd__mux2_1
X_5358_ _2084_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4309_ _2905_ _0386_ _2910_ _0390_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__o22ai_1
X_5289_ _2036_ _2034_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4660_ _1431_ _1433_ _1437_ _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3611_ BitStream_buffer.BitStream_buffer_valid_n vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4591_ _1370_ _1371_ _1372_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3542_ _2708_ _2601_ BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6261_ net63 _0276_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[38\] sky130_fd_sc_hd__dfxtp_2
X_3473_ _3006_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__clkbuf_2
X_6192_ net154 _0207_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[84\] sky130_fd_sc_hd__dfxtp_1
X_5212_ net10 _0770_ _1949_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__mux2_1
X_5143_ _0847_ _0343_ _0739_ _0346_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__o22ai_1
X_5074_ _2806_ _2752_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ _2707_ _2771_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4927_ BitStream_buffer.BS_buffer\[24\] _3047_ _3049_ BitStream_buffer.BS_buffer\[25\]
+ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _2723_ _2820_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__nand2_1
X_3809_ _2859_ BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4789_ _0514_ _2881_ _3024_ _2884_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2587_ _2587_ vssd1 vssd1 vccd1 vccd1 clknet_0__2587_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5830_ _2387_ _2383_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__nor2_1
X_5761_ _2381_ BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1 vccd1
+ _2386_ sky130_fd_sc_hd__nand2_1
X_4712_ _3060_ _3021_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__nor2_1
X_5692_ _2316_ _1102_ _1206_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4643_ _2757_ _2696_ _0440_ _2701_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4574_ _2856_ _3044_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3525_ _3053_ _3055_ _3056_ _3058_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6244_ net46 _0259_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[23\] sky130_fd_sc_hd__dfxtp_2
X_3456_ _2971_ _2978_ _2984_ _2989_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__or4_1
X_3387_ _2914_ _2916_ _2917_ _2920_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6175_ net137 _0190_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[101\] sky130_fd_sc_hd__dfxtp_2
X_5126_ _1900_ _1901_ _1902_ _1903_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__or4_1
X_5057_ _0560_ _2655_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__or2_1
X_4008_ BitStream_buffer.BS_buffer\[74\] _2679_ _2682_ BitStream_buffer.BS_buffer\[75\]
+ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__a22o_1
X_5959_ _2377_ _2373_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ _2794_ _2810_ _2826_ _2843_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ BitStream_buffer.BS_buffer\[66\] _3005_ BitStream_buffer.BS_buffer\[67\] _3008_
+ _1075_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__a221oi_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__inv_2
X_3172_ BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__clkbuf_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5813_ _2434_ _2436_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5744_ _2368_ _1934_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__nand2_1
X_5675_ _2117_ _1946_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4626_ _1402_ _1404_ _1406_ _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4557_ _2787_ BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__nand2_1
X_3508_ _2659_ _3020_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__and2_2
X_4488_ BitStream_buffer.BS_buffer\[52\] _2935_ BitStream_buffer.BS_buffer\[53\] _2938_
+ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a221oi_2
X_6227_ net189 _0242_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[49\] sky130_fd_sc_hd__dfxtp_4
X_3439_ _2659_ _2965_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__nand2_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ net120 _0173_ vssd1 vssd1 vccd1 vccd1 BitStream_buffer.BS_buffer\[118\] sky130_fd_sc_hd__dfxtp_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _0476_ _2889_ _1884_ _1885_ _1886_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 half_fill_counter[2] sky130_fd_sc_hd__buf_12
X_6093__24 clknet_1_1__leaf__2593_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__inv_2
X_6031__128 clknet_1_0__leaf__2587_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3790_ _2839_ _2784_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__or2_1
X_5994__94 clknet_1_0__leaf__2584_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5460_ _2153_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4411_ BitStream_buffer.BS_buffer\[27\] _0351_ BitStream_buffer.BS_buffer\[28\] _0354_
+ _1195_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__a221oi_1
X_5391_ _2108_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__inv_2
X_4342_ _2765_ _2714_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nand2_1
X_4273_ _0847_ _2916_ _0739_ _2920_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__o22ai_1
X_3224_ _2680_ _2711_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__nand2_2
.ends

