magic
tech sky130A
magscale 1 2
timestamp 1695390460
<< nwell >>
rect 1066 49221 48890 49542
rect 1066 48133 48890 48699
rect 1066 47045 48890 47611
rect 1066 45957 48890 46523
rect 1066 44869 48890 45435
rect 1066 43781 48890 44347
rect 1066 42693 48890 43259
rect 1066 41605 48890 42171
rect 1066 40517 48890 41083
rect 1066 39429 48890 39995
rect 1066 38341 48890 38907
rect 1066 37253 48890 37819
rect 1066 36165 48890 36731
rect 1066 35077 48890 35643
rect 1066 33989 48890 34555
rect 1066 32901 48890 33467
rect 1066 31813 48890 32379
rect 1066 30725 48890 31291
rect 1066 29637 48890 30203
rect 1066 28549 48890 29115
rect 1066 27461 48890 28027
rect 1066 26373 48890 26939
rect 1066 25285 48890 25851
rect 1066 24197 48890 24763
rect 1066 23109 48890 23675
rect 1066 22021 48890 22587
rect 1066 20933 48890 21499
rect 1066 19845 48890 20411
rect 1066 18757 48890 19323
rect 1066 17669 48890 18235
rect 1066 16581 48890 17147
rect 1066 15493 48890 16059
rect 1066 14405 48890 14971
rect 1066 13317 48890 13883
rect 1066 12229 48890 12795
rect 1066 11141 48890 11707
rect 1066 10053 48890 10619
rect 1066 8965 48890 9531
rect 1066 7877 48890 8443
rect 1066 6789 48890 7355
rect 1066 5701 48890 6267
rect 1066 4613 48890 5179
rect 1066 3525 48890 4091
rect 1066 2437 48890 3003
<< obsli1 >>
rect 1104 2159 48852 49521
<< obsm1 >>
rect 1104 1504 48852 49552
<< metal2 >>
rect 1490 0 1546 800
rect 2870 0 2926 800
rect 4250 0 4306 800
rect 5630 0 5686 800
rect 7010 0 7066 800
rect 8390 0 8446 800
rect 9770 0 9826 800
rect 11150 0 11206 800
rect 12530 0 12586 800
rect 13910 0 13966 800
rect 15290 0 15346 800
rect 16670 0 16726 800
rect 18050 0 18106 800
rect 19430 0 19486 800
rect 20810 0 20866 800
rect 22190 0 22246 800
rect 23570 0 23626 800
rect 24950 0 25006 800
rect 26330 0 26386 800
rect 27710 0 27766 800
rect 29090 0 29146 800
rect 30470 0 30526 800
rect 31850 0 31906 800
rect 33230 0 33286 800
rect 34610 0 34666 800
rect 35990 0 36046 800
rect 37370 0 37426 800
rect 38750 0 38806 800
rect 40130 0 40186 800
rect 41510 0 41566 800
rect 42890 0 42946 800
rect 44270 0 44326 800
rect 45650 0 45706 800
rect 47030 0 47086 800
rect 48410 0 48466 800
<< obsm2 >>
rect 1400 856 48452 49541
rect 1400 734 1434 856
rect 1602 734 2814 856
rect 2982 734 4194 856
rect 4362 734 5574 856
rect 5742 734 6954 856
rect 7122 734 8334 856
rect 8502 734 9714 856
rect 9882 734 11094 856
rect 11262 734 12474 856
rect 12642 734 13854 856
rect 14022 734 15234 856
rect 15402 734 16614 856
rect 16782 734 17994 856
rect 18162 734 19374 856
rect 19542 734 20754 856
rect 20922 734 22134 856
rect 22302 734 23514 856
rect 23682 734 24894 856
rect 25062 734 26274 856
rect 26442 734 27654 856
rect 27822 734 29034 856
rect 29202 734 30414 856
rect 30582 734 31794 856
rect 31962 734 33174 856
rect 33342 734 34554 856
rect 34722 734 35934 856
rect 36102 734 37314 856
rect 37482 734 38694 856
rect 38862 734 40074 856
rect 40242 734 41454 856
rect 41622 734 42834 856
rect 43002 734 44214 856
rect 44382 734 45594 856
rect 45762 734 46974 856
rect 47142 734 48354 856
<< obsm3 >>
rect 2497 1670 48379 49537
<< metal4 >>
rect 4208 2128 4528 49552
rect 19568 2128 19888 49552
rect 34928 2128 35248 49552
<< obsm4 >>
rect 3371 2211 4128 34645
rect 4608 2211 19488 34645
rect 19968 2211 34848 34645
rect 35328 2211 44101 34645
<< labels >>
rlabel metal2 s 4250 0 4306 800 6 BitStream_buffer_input[0]
port 1 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 BitStream_buffer_input[10]
port 2 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 BitStream_buffer_input[11]
port 3 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 BitStream_buffer_input[12]
port 4 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 BitStream_buffer_input[13]
port 5 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 BitStream_buffer_input[14]
port 6 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 BitStream_buffer_input[15]
port 7 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 BitStream_buffer_input[1]
port 8 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 BitStream_buffer_input[2]
port 9 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 BitStream_buffer_input[3]
port 10 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 BitStream_buffer_input[4]
port 11 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 BitStream_buffer_input[5]
port 12 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 BitStream_buffer_input[6]
port 13 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 BitStream_buffer_input[7]
port 14 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 BitStream_buffer_input[8]
port 15 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 BitStream_buffer_input[9]
port 16 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 clk
port 17 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 exp_golomb_decoding_output[0]
port 18 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 exp_golomb_decoding_output[1]
port 19 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 exp_golomb_decoding_output[2]
port 20 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 exp_golomb_decoding_output[3]
port 21 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 exp_golomb_decoding_output[4]
port 22 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 exp_golomb_decoding_output[5]
port 23 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 exp_golomb_decoding_output[6]
port 24 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 exp_golomb_decoding_output[7]
port 25 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 exp_golomb_sel[0]
port 26 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 exp_golomb_sel[1]
port 27 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 half_fill_counter[0]
port 28 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 half_fill_counter[1]
port 29 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 half_fill_counter[2]
port 30 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 reset_counter[0]
port 31 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 reset_counter[1]
port 32 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 reset_counter[2]
port 33 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 reset_counter[3]
port 34 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 reset_n
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 49552 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 49552 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 49552 6 vssd1
port 37 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 49973 52117
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9196374
string GDS_FILE /home/uniccass/H.264_Decoder/openlane/egd_top/runs/23_09_22_06_16/results/signoff/egd_top.magic.gds
string GDS_START 534066
<< end >>

