// This is the unpowered netlist.
module egd_top_wrapper (la_data_in_65,
    wb_clk_i,
    la_data_in_47_32,
    la_data_in_49_48,
    la_data_out_15_8,
    la_data_out_18_16,
    la_data_out_22_19);
 input la_data_in_65;
 input wb_clk_i;
 input [15:0] la_data_in_47_32;
 input [1:0] la_data_in_49_48;
 output [7:0] la_data_out_15_8;
 output [2:0] la_data_out_18_16;
 output [3:0] la_data_out_22_19;

 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire clknet_0__2958_;
 wire clknet_0__2959_;
 wire clknet_0__2960_;
 wire clknet_0__2961_;
 wire clknet_0__2962_;
 wire clknet_0__2963_;
 wire clknet_0__2964_;
 wire clknet_0__2965_;
 wire clknet_0__2966_;
 wire clknet_0__2967_;
 wire clknet_0__2968_;
 wire clknet_0__2969_;
 wire clknet_0__2970_;
 wire clknet_0__2971_;
 wire clknet_0__2972_;
 wire clknet_0__2973_;
 wire clknet_0__2974_;
 wire clknet_0__2975_;
 wire clknet_1_0__leaf__2958_;
 wire clknet_1_0__leaf__2959_;
 wire clknet_1_0__leaf__2960_;
 wire clknet_1_0__leaf__2961_;
 wire clknet_1_0__leaf__2962_;
 wire clknet_1_0__leaf__2963_;
 wire clknet_1_0__leaf__2964_;
 wire clknet_1_0__leaf__2965_;
 wire clknet_1_0__leaf__2966_;
 wire clknet_1_0__leaf__2967_;
 wire clknet_1_0__leaf__2968_;
 wire clknet_1_0__leaf__2969_;
 wire clknet_1_0__leaf__2970_;
 wire clknet_1_0__leaf__2971_;
 wire clknet_1_0__leaf__2972_;
 wire clknet_1_0__leaf__2973_;
 wire clknet_1_0__leaf__2974_;
 wire clknet_1_0__leaf__2975_;
 wire clknet_1_1__leaf__2958_;
 wire clknet_1_1__leaf__2959_;
 wire clknet_1_1__leaf__2960_;
 wire clknet_1_1__leaf__2961_;
 wire clknet_1_1__leaf__2962_;
 wire clknet_1_1__leaf__2963_;
 wire clknet_1_1__leaf__2964_;
 wire clknet_1_1__leaf__2965_;
 wire clknet_1_1__leaf__2966_;
 wire clknet_1_1__leaf__2967_;
 wire clknet_1_1__leaf__2968_;
 wire clknet_1_1__leaf__2969_;
 wire clknet_1_1__leaf__2970_;
 wire clknet_1_1__leaf__2971_;
 wire clknet_1_1__leaf__2972_;
 wire clknet_1_1__leaf__2973_;
 wire clknet_1_1__leaf__2974_;
 wire clknet_1_1__leaf__2975_;
 wire \egd_top.BitStream_buffer.BS_buffer[0] ;
 wire \egd_top.BitStream_buffer.BS_buffer[100] ;
 wire \egd_top.BitStream_buffer.BS_buffer[101] ;
 wire \egd_top.BitStream_buffer.BS_buffer[102] ;
 wire \egd_top.BitStream_buffer.BS_buffer[103] ;
 wire \egd_top.BitStream_buffer.BS_buffer[104] ;
 wire \egd_top.BitStream_buffer.BS_buffer[105] ;
 wire \egd_top.BitStream_buffer.BS_buffer[106] ;
 wire \egd_top.BitStream_buffer.BS_buffer[107] ;
 wire \egd_top.BitStream_buffer.BS_buffer[108] ;
 wire \egd_top.BitStream_buffer.BS_buffer[109] ;
 wire \egd_top.BitStream_buffer.BS_buffer[10] ;
 wire \egd_top.BitStream_buffer.BS_buffer[110] ;
 wire \egd_top.BitStream_buffer.BS_buffer[111] ;
 wire \egd_top.BitStream_buffer.BS_buffer[112] ;
 wire \egd_top.BitStream_buffer.BS_buffer[113] ;
 wire \egd_top.BitStream_buffer.BS_buffer[114] ;
 wire \egd_top.BitStream_buffer.BS_buffer[115] ;
 wire \egd_top.BitStream_buffer.BS_buffer[116] ;
 wire \egd_top.BitStream_buffer.BS_buffer[117] ;
 wire \egd_top.BitStream_buffer.BS_buffer[118] ;
 wire \egd_top.BitStream_buffer.BS_buffer[119] ;
 wire \egd_top.BitStream_buffer.BS_buffer[11] ;
 wire \egd_top.BitStream_buffer.BS_buffer[120] ;
 wire \egd_top.BitStream_buffer.BS_buffer[121] ;
 wire \egd_top.BitStream_buffer.BS_buffer[122] ;
 wire \egd_top.BitStream_buffer.BS_buffer[123] ;
 wire \egd_top.BitStream_buffer.BS_buffer[124] ;
 wire \egd_top.BitStream_buffer.BS_buffer[125] ;
 wire \egd_top.BitStream_buffer.BS_buffer[126] ;
 wire \egd_top.BitStream_buffer.BS_buffer[127] ;
 wire \egd_top.BitStream_buffer.BS_buffer[12] ;
 wire \egd_top.BitStream_buffer.BS_buffer[13] ;
 wire \egd_top.BitStream_buffer.BS_buffer[14] ;
 wire \egd_top.BitStream_buffer.BS_buffer[15] ;
 wire \egd_top.BitStream_buffer.BS_buffer[16] ;
 wire \egd_top.BitStream_buffer.BS_buffer[17] ;
 wire \egd_top.BitStream_buffer.BS_buffer[18] ;
 wire \egd_top.BitStream_buffer.BS_buffer[19] ;
 wire \egd_top.BitStream_buffer.BS_buffer[1] ;
 wire \egd_top.BitStream_buffer.BS_buffer[20] ;
 wire \egd_top.BitStream_buffer.BS_buffer[21] ;
 wire \egd_top.BitStream_buffer.BS_buffer[22] ;
 wire \egd_top.BitStream_buffer.BS_buffer[23] ;
 wire \egd_top.BitStream_buffer.BS_buffer[24] ;
 wire \egd_top.BitStream_buffer.BS_buffer[25] ;
 wire \egd_top.BitStream_buffer.BS_buffer[26] ;
 wire \egd_top.BitStream_buffer.BS_buffer[27] ;
 wire \egd_top.BitStream_buffer.BS_buffer[28] ;
 wire \egd_top.BitStream_buffer.BS_buffer[29] ;
 wire \egd_top.BitStream_buffer.BS_buffer[2] ;
 wire \egd_top.BitStream_buffer.BS_buffer[30] ;
 wire \egd_top.BitStream_buffer.BS_buffer[31] ;
 wire \egd_top.BitStream_buffer.BS_buffer[32] ;
 wire \egd_top.BitStream_buffer.BS_buffer[33] ;
 wire \egd_top.BitStream_buffer.BS_buffer[34] ;
 wire \egd_top.BitStream_buffer.BS_buffer[35] ;
 wire \egd_top.BitStream_buffer.BS_buffer[36] ;
 wire \egd_top.BitStream_buffer.BS_buffer[37] ;
 wire \egd_top.BitStream_buffer.BS_buffer[38] ;
 wire \egd_top.BitStream_buffer.BS_buffer[39] ;
 wire \egd_top.BitStream_buffer.BS_buffer[3] ;
 wire \egd_top.BitStream_buffer.BS_buffer[40] ;
 wire \egd_top.BitStream_buffer.BS_buffer[41] ;
 wire \egd_top.BitStream_buffer.BS_buffer[42] ;
 wire \egd_top.BitStream_buffer.BS_buffer[43] ;
 wire \egd_top.BitStream_buffer.BS_buffer[44] ;
 wire \egd_top.BitStream_buffer.BS_buffer[45] ;
 wire \egd_top.BitStream_buffer.BS_buffer[46] ;
 wire \egd_top.BitStream_buffer.BS_buffer[47] ;
 wire \egd_top.BitStream_buffer.BS_buffer[48] ;
 wire \egd_top.BitStream_buffer.BS_buffer[49] ;
 wire \egd_top.BitStream_buffer.BS_buffer[4] ;
 wire \egd_top.BitStream_buffer.BS_buffer[50] ;
 wire \egd_top.BitStream_buffer.BS_buffer[51] ;
 wire \egd_top.BitStream_buffer.BS_buffer[52] ;
 wire \egd_top.BitStream_buffer.BS_buffer[53] ;
 wire \egd_top.BitStream_buffer.BS_buffer[54] ;
 wire \egd_top.BitStream_buffer.BS_buffer[55] ;
 wire \egd_top.BitStream_buffer.BS_buffer[56] ;
 wire \egd_top.BitStream_buffer.BS_buffer[57] ;
 wire \egd_top.BitStream_buffer.BS_buffer[58] ;
 wire \egd_top.BitStream_buffer.BS_buffer[59] ;
 wire \egd_top.BitStream_buffer.BS_buffer[5] ;
 wire \egd_top.BitStream_buffer.BS_buffer[60] ;
 wire \egd_top.BitStream_buffer.BS_buffer[61] ;
 wire \egd_top.BitStream_buffer.BS_buffer[62] ;
 wire \egd_top.BitStream_buffer.BS_buffer[63] ;
 wire \egd_top.BitStream_buffer.BS_buffer[64] ;
 wire \egd_top.BitStream_buffer.BS_buffer[65] ;
 wire \egd_top.BitStream_buffer.BS_buffer[66] ;
 wire \egd_top.BitStream_buffer.BS_buffer[67] ;
 wire \egd_top.BitStream_buffer.BS_buffer[68] ;
 wire \egd_top.BitStream_buffer.BS_buffer[69] ;
 wire \egd_top.BitStream_buffer.BS_buffer[6] ;
 wire \egd_top.BitStream_buffer.BS_buffer[70] ;
 wire \egd_top.BitStream_buffer.BS_buffer[71] ;
 wire \egd_top.BitStream_buffer.BS_buffer[72] ;
 wire \egd_top.BitStream_buffer.BS_buffer[73] ;
 wire \egd_top.BitStream_buffer.BS_buffer[74] ;
 wire \egd_top.BitStream_buffer.BS_buffer[75] ;
 wire \egd_top.BitStream_buffer.BS_buffer[76] ;
 wire \egd_top.BitStream_buffer.BS_buffer[77] ;
 wire \egd_top.BitStream_buffer.BS_buffer[78] ;
 wire \egd_top.BitStream_buffer.BS_buffer[79] ;
 wire \egd_top.BitStream_buffer.BS_buffer[7] ;
 wire \egd_top.BitStream_buffer.BS_buffer[80] ;
 wire \egd_top.BitStream_buffer.BS_buffer[81] ;
 wire \egd_top.BitStream_buffer.BS_buffer[82] ;
 wire \egd_top.BitStream_buffer.BS_buffer[83] ;
 wire \egd_top.BitStream_buffer.BS_buffer[84] ;
 wire \egd_top.BitStream_buffer.BS_buffer[85] ;
 wire \egd_top.BitStream_buffer.BS_buffer[86] ;
 wire \egd_top.BitStream_buffer.BS_buffer[87] ;
 wire \egd_top.BitStream_buffer.BS_buffer[88] ;
 wire \egd_top.BitStream_buffer.BS_buffer[89] ;
 wire \egd_top.BitStream_buffer.BS_buffer[8] ;
 wire \egd_top.BitStream_buffer.BS_buffer[90] ;
 wire \egd_top.BitStream_buffer.BS_buffer[91] ;
 wire \egd_top.BitStream_buffer.BS_buffer[92] ;
 wire \egd_top.BitStream_buffer.BS_buffer[93] ;
 wire \egd_top.BitStream_buffer.BS_buffer[94] ;
 wire \egd_top.BitStream_buffer.BS_buffer[95] ;
 wire \egd_top.BitStream_buffer.BS_buffer[96] ;
 wire \egd_top.BitStream_buffer.BS_buffer[97] ;
 wire \egd_top.BitStream_buffer.BS_buffer[98] ;
 wire \egd_top.BitStream_buffer.BS_buffer[99] ;
 wire \egd_top.BitStream_buffer.BS_buffer[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[10] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[11] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[12] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[13] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[14] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[15] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[1] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[2] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[3] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[4] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[5] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[6] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[7] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[8] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_valid_n ;
 wire \egd_top.BitStream_buffer.buffer_index[4] ;
 wire \egd_top.BitStream_buffer.buffer_index[5] ;
 wire \egd_top.BitStream_buffer.buffer_index[6] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[1] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[2] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[3] ;
 wire \egd_top.BitStream_buffer.pc[1] ;
 wire \egd_top.BitStream_buffer.pc[2] ;
 wire \egd_top.BitStream_buffer.pc[3] ;
 wire \egd_top.BitStream_buffer.pc[4] ;
 wire \egd_top.BitStream_buffer.pc[5] ;
 wire \egd_top.BitStream_buffer.pc[6] ;
 wire \egd_top.BitStream_buffer.pc_previous[0] ;
 wire \egd_top.BitStream_buffer.pc_previous[1] ;
 wire \egd_top.BitStream_buffer.pc_previous[2] ;
 wire \egd_top.BitStream_buffer.pc_previous[3] ;
 wire \egd_top.BitStream_buffer.pc_previous[4] ;
 wire \egd_top.BitStream_buffer.pc_previous[5] ;
 wire \egd_top.BitStream_buffer.pc_previous[6] ;
 wire \egd_top.exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net14));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_92 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__inv_2 _3418_ (.A(net33),
    .Y(_2976_));
 sky130_fd_sc_hd__nand2_1 _3419_ (.A(net32),
    .B(net31),
    .Y(_2977_));
 sky130_fd_sc_hd__inv_2 _3420_ (.A(net34),
    .Y(_2978_));
 sky130_fd_sc_hd__o21ai_1 _3421_ (.A1(_2976_),
    .A2(_2977_),
    .B1(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__buf_2 _3422_ (.A(net19),
    .X(_2980_));
 sky130_fd_sc_hd__and2_1 _3423_ (.A(_2979_),
    .B(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__clkbuf_1 _3424_ (.A(_2981_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _3425_ (.A1(_2976_),
    .A2(_2977_),
    .B1(_2979_),
    .X(_2982_));
 sky130_fd_sc_hd__nand2_1 _3426_ (.A(net34),
    .B(net33),
    .Y(_2983_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(net19),
    .Y(_2984_));
 sky130_fd_sc_hd__clkbuf_4 _3428_ (.A(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__a21oi_1 _3429_ (.A1(_2982_),
    .A2(_2983_),
    .B1(_2985_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _3430_ (.A(net31),
    .Y(_2986_));
 sky130_fd_sc_hd__nor2_1 _3431_ (.A(net33),
    .B(net32),
    .Y(_2987_));
 sky130_fd_sc_hd__nor2_1 _3432_ (.A(_2978_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__nor2_1 _3433_ (.A(_2986_),
    .B(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__a21o_1 _3434_ (.A1(_2989_),
    .A2(net32),
    .B1(_2984_),
    .X(_2990_));
 sky130_fd_sc_hd__o21ba_1 _3435_ (.A1(net32),
    .A2(_2989_),
    .B1_N(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__clkbuf_1 _3436_ (.A(_2991_),
    .X(_0319_));
 sky130_fd_sc_hd__inv_2 _3437_ (.A(_2988_),
    .Y(_2992_));
 sky130_fd_sc_hd__nor2_1 _3438_ (.A(net31),
    .B(_2992_),
    .Y(_2993_));
 sky130_fd_sc_hd__or3_1 _3439_ (.A(_2984_),
    .B(_2989_),
    .C(_2993_),
    .X(_2994_));
 sky130_fd_sc_hd__inv_2 _3440_ (.A(_2994_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _3441_ (.A(net30),
    .Y(_2995_));
 sky130_fd_sc_hd__nor2_1 _3442_ (.A(net29),
    .B(net28),
    .Y(_2996_));
 sky130_fd_sc_hd__nor2_1 _3443_ (.A(_2995_),
    .B(_2996_),
    .Y(_2997_));
 sky130_fd_sc_hd__a21o_1 _3444_ (.A1(net29),
    .A2(net28),
    .B1(net30),
    .X(_2998_));
 sky130_fd_sc_hd__and2b_1 _3445_ (.A_N(_2997_),
    .B(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__inv_2 _3446_ (.A(net29),
    .Y(_3000_));
 sky130_fd_sc_hd__nand2_4 _3447_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3001_));
 sky130_fd_sc_hd__inv_2 _3448_ (.A(net18),
    .Y(_3002_));
 sky130_fd_sc_hd__inv_4 _3449_ (.A(net17),
    .Y(_3003_));
 sky130_fd_sc_hd__nand2_2 _3450_ (.A(_3002_),
    .B(_3003_),
    .Y(_3004_));
 sky130_fd_sc_hd__or2_1 _3451_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__nand2_4 _3452_ (.A(_3004_),
    .B(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_3006_));
 sky130_fd_sc_hd__nand2_2 _3453_ (.A(_3005_),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__inv_2 _3454_ (.A(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__nand2_2 _3455_ (.A(_3008_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3009_));
 sky130_fd_sc_hd__nor2_4 _3456_ (.A(_3001_),
    .B(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__inv_2 _3457_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_3011_));
 sky130_fd_sc_hd__and3_1 _3458_ (.A(_3011_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3012_));
 sky130_fd_sc_hd__and2_1 _3459_ (.A(_3010_),
    .B(_3012_),
    .X(_3013_));
 sky130_fd_sc_hd__nor2_1 _3460_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_3013_),
    .Y(_3014_));
 sky130_fd_sc_hd__inv_2 _3461_ (.A(_2996_),
    .Y(_3015_));
 sky130_fd_sc_hd__nor2_1 _3462_ (.A(net30),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__inv_2 _3463_ (.A(net198),
    .Y(_3017_));
 sky130_fd_sc_hd__inv_2 _3464_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_3018_));
 sky130_fd_sc_hd__and3_1 _3465_ (.A(_3017_),
    .B(_3018_),
    .C(net196),
    .X(_3019_));
 sky130_fd_sc_hd__nand3_1 _3466_ (.A(_3014_),
    .B(_3016_),
    .C(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__nor2_1 _3467_ (.A(_2997_),
    .B(_3016_),
    .Y(_3021_));
 sky130_fd_sc_hd__inv_2 _3468_ (.A(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__nand2_1 _3469_ (.A(_3020_),
    .B(_3022_),
    .Y(_3023_));
 sky130_fd_sc_hd__inv_2 _3470_ (.A(net196),
    .Y(_3024_));
 sky130_fd_sc_hd__and3_1 _3471_ (.A(_3024_),
    .B(_3017_),
    .C(_3018_),
    .X(_3025_));
 sky130_fd_sc_hd__and4_1 _3472_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(\egd_top.BitStream_buffer.pc_previous[1] ),
    .C(\egd_top.BitStream_buffer.pc_previous[2] ),
    .D(\egd_top.BitStream_buffer.pc_previous[3] ),
    .X(_3026_));
 sky130_fd_sc_hd__a31o_1 _3473_ (.A1(_3026_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .A3(\egd_top.BitStream_buffer.pc_previous[5] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[6] ),
    .X(_3027_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(_3014_),
    .B(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__or2_1 _3475_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_3011_),
    .X(_3029_));
 sky130_fd_sc_hd__a21boi_1 _3476_ (.A1(_3028_),
    .A2(_3029_),
    .B1_N(_3016_),
    .Y(_3030_));
 sky130_fd_sc_hd__a31o_1 _3477_ (.A1(\egd_top.BitStream_buffer.pc[6] ),
    .A2(_3016_),
    .A3(_3025_),
    .B1(_3030_),
    .X(_3031_));
 sky130_fd_sc_hd__a311o_1 _3478_ (.A1(net30),
    .A2(_3000_),
    .A3(net28),
    .B1(_3023_),
    .C1(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__and4_1 _3479_ (.A(_2976_),
    .B(_2986_),
    .C(net34),
    .D(net32),
    .X(_3033_));
 sky130_fd_sc_hd__nand2_2 _3480_ (.A(_3032_),
    .B(_3033_),
    .Y(_3034_));
 sky130_fd_sc_hd__buf_4 _3481_ (.A(net19),
    .X(_3035_));
 sky130_fd_sc_hd__buf_2 _3482_ (.A(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__nand2_1 _3483_ (.A(_3034_),
    .B(_2995_),
    .Y(_3037_));
 sky130_fd_sc_hd__o211a_1 _3484_ (.A1(_2999_),
    .A2(_3034_),
    .B1(_3036_),
    .C1(_3037_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _3485_ (.A(_2996_),
    .B(_2998_),
    .Y(_3038_));
 sky130_fd_sc_hd__nand2_1 _3486_ (.A(_3034_),
    .B(_3000_),
    .Y(_3039_));
 sky130_fd_sc_hd__o211a_1 _3487_ (.A1(_3038_),
    .A2(_3034_),
    .B1(_3036_),
    .C1(_3039_),
    .X(_0316_));
 sky130_fd_sc_hd__o21ai_1 _3488_ (.A1(net28),
    .A2(_3022_),
    .B1(_3020_),
    .Y(_3040_));
 sky130_fd_sc_hd__o21bai_1 _3489_ (.A1(_3031_),
    .A2(_3040_),
    .B1_N(_3034_),
    .Y(_3041_));
 sky130_fd_sc_hd__nand2_1 _3490_ (.A(_3034_),
    .B(net28),
    .Y(_3042_));
 sky130_fd_sc_hd__a21oi_1 _3491_ (.A1(_3041_),
    .A2(_3042_),
    .B1(_2985_),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _3492_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .Y(_3043_));
 sky130_fd_sc_hd__o21ai_1 _3493_ (.A1(_3043_),
    .A2(_3033_),
    .B1(_3036_),
    .Y(_0314_));
 sky130_fd_sc_hd__buf_2 _3494_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .X(_3044_));
 sky130_fd_sc_hd__nand2_1 _3495_ (.A(_2995_),
    .B(_3000_),
    .Y(_3045_));
 sky130_fd_sc_hd__nand2_1 _3496_ (.A(net30),
    .B(net202),
    .Y(_3046_));
 sky130_fd_sc_hd__nand2_1 _3497_ (.A(_2987_),
    .B(_2978_),
    .Y(_3047_));
 sky130_fd_sc_hd__a22o_4 _3498_ (.A1(_3045_),
    .A2(_3046_),
    .B1(_2992_),
    .B2(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__nand2_1 _3499_ (.A(_3048_),
    .B(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_3049_));
 sky130_fd_sc_hd__or2_1 _3500_ (.A(_3017_),
    .B(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__or2_1 _3501_ (.A(_3024_),
    .B(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__buf_2 _3502_ (.A(_3051_),
    .X(_3052_));
 sky130_fd_sc_hd__clkbuf_4 _3503_ (.A(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(net7),
    .A1(_3044_),
    .S(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__and2_1 _3505_ (.A(_3054_),
    .B(_2980_),
    .X(_3055_));
 sky130_fd_sc_hd__clkbuf_1 _3506_ (.A(_3055_),
    .X(_0313_));
 sky130_fd_sc_hd__buf_2 _3507_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_3056_));
 sky130_fd_sc_hd__mux2_1 _3508_ (.A0(net6),
    .A1(_3056_),
    .S(_3053_),
    .X(_3057_));
 sky130_fd_sc_hd__and2_1 _3509_ (.A(_3057_),
    .B(_2980_),
    .X(_3058_));
 sky130_fd_sc_hd__clkbuf_1 _3510_ (.A(_3058_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_2 _3511_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .X(_3059_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(net5),
    .A1(_3059_),
    .S(_3053_),
    .X(_3060_));
 sky130_fd_sc_hd__and2_1 _3513_ (.A(_3060_),
    .B(_2980_),
    .X(_3061_));
 sky130_fd_sc_hd__clkbuf_1 _3514_ (.A(_3061_),
    .X(_0311_));
 sky130_fd_sc_hd__buf_2 _3515_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .X(_3062_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(net4),
    .A1(_3062_),
    .S(_3053_),
    .X(_3063_));
 sky130_fd_sc_hd__and2_1 _3517_ (.A(_3063_),
    .B(_2980_),
    .X(_3064_));
 sky130_fd_sc_hd__clkbuf_1 _3518_ (.A(_3064_),
    .X(_0310_));
 sky130_fd_sc_hd__buf_2 _3519_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .X(_3065_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(net3),
    .A1(_3065_),
    .S(_3053_),
    .X(_3066_));
 sky130_fd_sc_hd__and2_1 _3521_ (.A(_3066_),
    .B(_2980_),
    .X(_3067_));
 sky130_fd_sc_hd__clkbuf_1 _3522_ (.A(_3067_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_2 _3523_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .X(_3068_));
 sky130_fd_sc_hd__mux2_1 _3524_ (.A0(net2),
    .A1(_3068_),
    .S(_3053_),
    .X(_3069_));
 sky130_fd_sc_hd__and2_1 _3525_ (.A(_3069_),
    .B(_2980_),
    .X(_3070_));
 sky130_fd_sc_hd__clkbuf_1 _3526_ (.A(_3070_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_4 _3527_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .X(_3071_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(net16),
    .A1(_3071_),
    .S(_3053_),
    .X(_3072_));
 sky130_fd_sc_hd__and2_1 _3529_ (.A(_3072_),
    .B(_2980_),
    .X(_3073_));
 sky130_fd_sc_hd__clkbuf_1 _3530_ (.A(_3073_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_2 _3531_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_3074_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(net15),
    .A1(_3074_),
    .S(_3053_),
    .X(_3075_));
 sky130_fd_sc_hd__clkbuf_2 _3533_ (.A(_3035_),
    .X(_3076_));
 sky130_fd_sc_hd__and2_1 _3534_ (.A(_3075_),
    .B(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__clkbuf_1 _3535_ (.A(_3077_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_2 _3536_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_3078_));
 sky130_fd_sc_hd__mux2_1 _3537_ (.A0(net14),
    .A1(_3078_),
    .S(_3053_),
    .X(_3079_));
 sky130_fd_sc_hd__and2_1 _3538_ (.A(_3079_),
    .B(_3076_),
    .X(_3080_));
 sky130_fd_sc_hd__clkbuf_1 _3539_ (.A(_3080_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_2 _3540_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_3081_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(net13),
    .A1(_3081_),
    .S(_3052_),
    .X(_3082_));
 sky130_fd_sc_hd__and2_1 _3542_ (.A(_3082_),
    .B(_3076_),
    .X(_3083_));
 sky130_fd_sc_hd__clkbuf_1 _3543_ (.A(_3083_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_4 _3544_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_3084_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(net12),
    .A1(_3084_),
    .S(_3052_),
    .X(_3085_));
 sky130_fd_sc_hd__and2_1 _3546_ (.A(_3085_),
    .B(_3076_),
    .X(_3086_));
 sky130_fd_sc_hd__clkbuf_1 _3547_ (.A(_3086_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_4 _3548_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .X(_3087_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(net11),
    .A1(_3087_),
    .S(_3052_),
    .X(_3088_));
 sky130_fd_sc_hd__and2_1 _3550_ (.A(_3088_),
    .B(_3076_),
    .X(_3089_));
 sky130_fd_sc_hd__clkbuf_1 _3551_ (.A(_3089_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_2 _3552_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_3090_));
 sky130_fd_sc_hd__mux2_1 _3553_ (.A0(net10),
    .A1(_3090_),
    .S(_3052_),
    .X(_3091_));
 sky130_fd_sc_hd__and2_1 _3554_ (.A(_3091_),
    .B(_3076_),
    .X(_3092_));
 sky130_fd_sc_hd__clkbuf_1 _3555_ (.A(_3092_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_4 _3556_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_3093_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(net9),
    .A1(_3093_),
    .S(_3052_),
    .X(_3094_));
 sky130_fd_sc_hd__and2_1 _3558_ (.A(_3094_),
    .B(_3076_),
    .X(_3095_));
 sky130_fd_sc_hd__clkbuf_1 _3559_ (.A(_3095_),
    .X(_0300_));
 sky130_fd_sc_hd__buf_2 _3560_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_3096_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(net8),
    .A1(_3096_),
    .S(_3052_),
    .X(_3097_));
 sky130_fd_sc_hd__and2_1 _3562_ (.A(_3097_),
    .B(_3076_),
    .X(_3098_));
 sky130_fd_sc_hd__clkbuf_1 _3563_ (.A(_3098_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_2 _3564_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_3099_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(net1),
    .A1(_3099_),
    .S(_3052_),
    .X(_3100_));
 sky130_fd_sc_hd__and2_1 _3566_ (.A(_3100_),
    .B(_3076_),
    .X(_3101_));
 sky130_fd_sc_hd__clkbuf_1 _3567_ (.A(_3101_),
    .X(_0298_));
 sky130_fd_sc_hd__buf_2 _3568_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .X(_3102_));
 sky130_fd_sc_hd__buf_2 _3569_ (.A(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__buf_2 _3570_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_3104_));
 sky130_fd_sc_hd__nand2_2 _3571_ (.A(_3007_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3105_));
 sky130_fd_sc_hd__inv_2 _3572_ (.A(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__inv_2 _3573_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_3107_));
 sky130_fd_sc_hd__and3_2 _3574_ (.A(_3106_),
    .B(_3107_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3108_));
 sky130_fd_sc_hd__inv_2 _3575_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_3109_));
 sky130_fd_sc_hd__inv_2 _3576_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_3110_));
 sky130_fd_sc_hd__and3_1 _3577_ (.A(_3109_),
    .B(_3110_),
    .C(\egd_top.BitStream_buffer.pc[6] ),
    .X(_3111_));
 sky130_fd_sc_hd__clkbuf_4 _3578_ (.A(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__and2_1 _3579_ (.A(_3108_),
    .B(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__clkbuf_2 _3580_ (.A(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__buf_2 _3581_ (.A(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__buf_2 _3582_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_3116_));
 sky130_fd_sc_hd__inv_2 _3583_ (.A(_3009_),
    .Y(_3117_));
 sky130_fd_sc_hd__and3_1 _3584_ (.A(_3117_),
    .B(_3107_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3118_));
 sky130_fd_sc_hd__buf_6 _3585_ (.A(_3118_),
    .X(_3119_));
 sky130_fd_sc_hd__and2_1 _3586_ (.A(_3119_),
    .B(_3112_),
    .X(_3120_));
 sky130_fd_sc_hd__clkbuf_2 _3587_ (.A(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__buf_4 _3588_ (.A(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__inv_2 _3589_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_3123_));
 sky130_fd_sc_hd__inv_2 _3590_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3124_));
 sky130_fd_sc_hd__nand2_2 _3591_ (.A(_3007_),
    .B(_3124_),
    .Y(_3125_));
 sky130_fd_sc_hd__inv_2 _3592_ (.A(_3125_),
    .Y(_3126_));
 sky130_fd_sc_hd__and3_1 _3593_ (.A(_3126_),
    .B(_3107_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3127_));
 sky130_fd_sc_hd__buf_4 _3594_ (.A(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__nand2_2 _3595_ (.A(_3128_),
    .B(_3112_),
    .Y(_3129_));
 sky130_fd_sc_hd__buf_2 _3596_ (.A(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__clkbuf_4 _3597_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_3131_));
 sky130_fd_sc_hd__inv_2 _3598_ (.A(_3131_),
    .Y(_3132_));
 sky130_fd_sc_hd__nand2_2 _3599_ (.A(_3008_),
    .B(_3124_),
    .Y(_3133_));
 sky130_fd_sc_hd__inv_2 _3600_ (.A(_3133_),
    .Y(_3134_));
 sky130_fd_sc_hd__and3_1 _3601_ (.A(_3134_),
    .B(_3107_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3135_));
 sky130_fd_sc_hd__clkbuf_4 _3602_ (.A(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__nand2_2 _3603_ (.A(_3136_),
    .B(_3112_),
    .Y(_3137_));
 sky130_fd_sc_hd__buf_2 _3604_ (.A(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__o22ai_1 _3605_ (.A1(_3123_),
    .A2(_3130_),
    .B1(_3132_),
    .B2(_3138_),
    .Y(_3139_));
 sky130_fd_sc_hd__a221oi_1 _3606_ (.A1(_3104_),
    .A2(_3115_),
    .B1(_3116_),
    .B2(_3122_),
    .C1(_3139_),
    .Y(_3140_));
 sky130_fd_sc_hd__buf_2 _3607_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .X(_3141_));
 sky130_fd_sc_hd__inv_2 _3608_ (.A(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3142_));
 sky130_fd_sc_hd__nand2_4 _3609_ (.A(_3107_),
    .B(_3142_),
    .Y(_3143_));
 sky130_fd_sc_hd__nor2_4 _3610_ (.A(_3143_),
    .B(_3105_),
    .Y(_3144_));
 sky130_fd_sc_hd__and2_1 _3611_ (.A(_3144_),
    .B(_3112_),
    .X(_3145_));
 sky130_fd_sc_hd__clkbuf_2 _3612_ (.A(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__buf_2 _3613_ (.A(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__buf_2 _3614_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .X(_3148_));
 sky130_fd_sc_hd__nor2_2 _3615_ (.A(_3143_),
    .B(_3009_),
    .Y(_3149_));
 sky130_fd_sc_hd__and2_1 _3616_ (.A(_3149_),
    .B(_3112_),
    .X(_3150_));
 sky130_fd_sc_hd__clkbuf_2 _3617_ (.A(_3150_),
    .X(_3151_));
 sky130_fd_sc_hd__clkbuf_4 _3618_ (.A(_3151_),
    .X(_3152_));
 sky130_fd_sc_hd__inv_2 _3619_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_3153_));
 sky130_fd_sc_hd__nor2_4 _3620_ (.A(_3143_),
    .B(_3125_),
    .Y(_3154_));
 sky130_fd_sc_hd__nand2_2 _3621_ (.A(_3154_),
    .B(_3112_),
    .Y(_3155_));
 sky130_fd_sc_hd__buf_2 _3622_ (.A(_3155_),
    .X(_3156_));
 sky130_fd_sc_hd__nor2_4 _3623_ (.A(_3143_),
    .B(_3133_),
    .Y(_3157_));
 sky130_fd_sc_hd__and2_1 _3624_ (.A(_3157_),
    .B(_3111_),
    .X(_3158_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3625_ (.A(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__buf_2 _3626_ (.A(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__buf_2 _3627_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .X(_3161_));
 sky130_fd_sc_hd__nand2_1 _3628_ (.A(_3160_),
    .B(_3161_),
    .Y(_3162_));
 sky130_fd_sc_hd__o21ai_1 _3629_ (.A1(_3153_),
    .A2(_3156_),
    .B1(_3162_),
    .Y(_3163_));
 sky130_fd_sc_hd__a221oi_1 _3630_ (.A1(_3141_),
    .A2(_3147_),
    .B1(_3148_),
    .B2(_3152_),
    .C1(_3163_),
    .Y(_3164_));
 sky130_fd_sc_hd__inv_2 _3631_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_3165_));
 sky130_fd_sc_hd__and3_1 _3632_ (.A(_3117_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3142_),
    .X(_3166_));
 sky130_fd_sc_hd__clkbuf_4 _3633_ (.A(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__nand2_2 _3634_ (.A(_3167_),
    .B(_3112_),
    .Y(_3168_));
 sky130_fd_sc_hd__buf_2 _3635_ (.A(_3168_),
    .X(_3169_));
 sky130_fd_sc_hd__and3_1 _3636_ (.A(_3126_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3142_),
    .X(_3170_));
 sky130_fd_sc_hd__clkbuf_4 _3637_ (.A(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__and2_1 _3638_ (.A(_3171_),
    .B(_3111_),
    .X(_3172_));
 sky130_fd_sc_hd__clkbuf_2 _3639_ (.A(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__buf_2 _3640_ (.A(_3173_),
    .X(_3174_));
 sky130_fd_sc_hd__buf_2 _3641_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .X(_3175_));
 sky130_fd_sc_hd__nand2_1 _3642_ (.A(_3174_),
    .B(_3175_),
    .Y(_3176_));
 sky130_fd_sc_hd__and3_2 _3643_ (.A(_3106_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3142_),
    .X(_3177_));
 sky130_fd_sc_hd__and2_1 _3644_ (.A(_3177_),
    .B(_3111_),
    .X(_3178_));
 sky130_fd_sc_hd__clkbuf_2 _3645_ (.A(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__buf_2 _3646_ (.A(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__buf_2 _3647_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_3181_));
 sky130_fd_sc_hd__nand2_1 _3648_ (.A(_3180_),
    .B(_3181_),
    .Y(_3182_));
 sky130_fd_sc_hd__inv_2 _3649_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_3183_));
 sky130_fd_sc_hd__and3_1 _3650_ (.A(_3134_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3142_),
    .X(_3184_));
 sky130_fd_sc_hd__buf_4 _3651_ (.A(_3184_),
    .X(_3185_));
 sky130_fd_sc_hd__nand2_2 _3652_ (.A(_3185_),
    .B(_3112_),
    .Y(_3186_));
 sky130_fd_sc_hd__clkbuf_2 _3653_ (.A(_3186_),
    .X(_3187_));
 sky130_fd_sc_hd__or2_1 _3654_ (.A(_3183_),
    .B(_3187_),
    .X(_3188_));
 sky130_fd_sc_hd__o2111a_1 _3655_ (.A1(_3165_),
    .A2(_3169_),
    .B1(_3176_),
    .C1(_3182_),
    .D1(_3188_),
    .X(_3189_));
 sky130_fd_sc_hd__buf_2 _3656_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_3190_));
 sky130_fd_sc_hd__nor2_4 _3657_ (.A(_3001_),
    .B(_3105_),
    .Y(_3191_));
 sky130_fd_sc_hd__and2_1 _3658_ (.A(_3191_),
    .B(_3111_),
    .X(_3192_));
 sky130_fd_sc_hd__clkbuf_2 _3659_ (.A(_3192_),
    .X(_3193_));
 sky130_fd_sc_hd__buf_4 _3660_ (.A(_3193_),
    .X(_3194_));
 sky130_fd_sc_hd__buf_2 _3661_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_3195_));
 sky130_fd_sc_hd__and2_1 _3662_ (.A(_3010_),
    .B(_3112_),
    .X(_3196_));
 sky130_fd_sc_hd__clkbuf_2 _3663_ (.A(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__buf_4 _3664_ (.A(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__nor2_4 _3665_ (.A(_3001_),
    .B(_3133_),
    .Y(_3199_));
 sky130_fd_sc_hd__and2_1 _3666_ (.A(_3199_),
    .B(_3111_),
    .X(_3200_));
 sky130_fd_sc_hd__clkbuf_2 _3667_ (.A(_3200_),
    .X(_3201_));
 sky130_fd_sc_hd__buf_2 _3668_ (.A(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__clkbuf_4 _3669_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_3203_));
 sky130_fd_sc_hd__nand2_1 _3670_ (.A(_3202_),
    .B(_3203_),
    .Y(_3204_));
 sky130_fd_sc_hd__nor2_4 _3671_ (.A(_3001_),
    .B(_3125_),
    .Y(_3205_));
 sky130_fd_sc_hd__and2_1 _3672_ (.A(_3205_),
    .B(_3111_),
    .X(_3206_));
 sky130_fd_sc_hd__clkbuf_2 _3673_ (.A(_3206_),
    .X(_3207_));
 sky130_fd_sc_hd__buf_2 _3674_ (.A(_3207_),
    .X(_3208_));
 sky130_fd_sc_hd__clkbuf_4 _3675_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_3209_));
 sky130_fd_sc_hd__nand2_1 _3676_ (.A(_3208_),
    .B(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__nand2_1 _3677_ (.A(_3204_),
    .B(_3210_),
    .Y(_3211_));
 sky130_fd_sc_hd__a221oi_1 _3678_ (.A1(_3190_),
    .A2(_3194_),
    .B1(_3195_),
    .B2(_3198_),
    .C1(_3211_),
    .Y(_3212_));
 sky130_fd_sc_hd__and4_1 _3679_ (.A(_3140_),
    .B(_3164_),
    .C(_3189_),
    .D(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__and3_2 _3680_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3214_));
 sky130_fd_sc_hd__clkbuf_4 _3681_ (.A(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__and2_1 _3682_ (.A(_3177_),
    .B(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__clkbuf_2 _3683_ (.A(_3216_),
    .X(_3217_));
 sky130_fd_sc_hd__buf_2 _3684_ (.A(_3217_),
    .X(_3218_));
 sky130_fd_sc_hd__and2_1 _3685_ (.A(_3167_),
    .B(_3215_),
    .X(_3219_));
 sky130_fd_sc_hd__clkbuf_2 _3686_ (.A(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__buf_6 _3687_ (.A(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__inv_2 _3688_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_3222_));
 sky130_fd_sc_hd__nand2_2 _3689_ (.A(_3171_),
    .B(_3215_),
    .Y(_3223_));
 sky130_fd_sc_hd__buf_2 _3690_ (.A(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__inv_2 _3691_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_3225_));
 sky130_fd_sc_hd__nand2_2 _3692_ (.A(_3185_),
    .B(_3215_),
    .Y(_3226_));
 sky130_fd_sc_hd__buf_2 _3693_ (.A(_3226_),
    .X(_3227_));
 sky130_fd_sc_hd__o22ai_1 _3694_ (.A1(_3222_),
    .A2(_3224_),
    .B1(_3225_),
    .B2(_3227_),
    .Y(_3228_));
 sky130_fd_sc_hd__a221oi_1 _3695_ (.A1(_3071_),
    .A2(_3218_),
    .B1(_3074_),
    .B2(_3221_),
    .C1(_3228_),
    .Y(_3229_));
 sky130_fd_sc_hd__and2_1 _3696_ (.A(_3128_),
    .B(_3214_),
    .X(_3230_));
 sky130_fd_sc_hd__clkbuf_2 _3697_ (.A(_3230_),
    .X(_3231_));
 sky130_fd_sc_hd__clkbuf_4 _3698_ (.A(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__and2_1 _3699_ (.A(_3136_),
    .B(_3215_),
    .X(_3233_));
 sky130_fd_sc_hd__clkbuf_2 _3700_ (.A(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__buf_4 _3701_ (.A(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__inv_2 _3702_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_3236_));
 sky130_fd_sc_hd__nand2_2 _3703_ (.A(_3119_),
    .B(_3215_),
    .Y(_3237_));
 sky130_fd_sc_hd__clkbuf_4 _3704_ (.A(_3237_),
    .X(_3238_));
 sky130_fd_sc_hd__and2_1 _3705_ (.A(_3108_),
    .B(_3214_),
    .X(_3239_));
 sky130_fd_sc_hd__clkbuf_2 _3706_ (.A(_3239_),
    .X(_3240_));
 sky130_fd_sc_hd__buf_2 _3707_ (.A(_3240_),
    .X(_3241_));
 sky130_fd_sc_hd__nand2_1 _3708_ (.A(_3241_),
    .B(_3084_),
    .Y(_3242_));
 sky130_fd_sc_hd__o21ai_1 _3709_ (.A1(_3236_),
    .A2(_3238_),
    .B1(_3242_),
    .Y(_3243_));
 sky130_fd_sc_hd__a221oi_1 _3710_ (.A1(_3078_),
    .A2(_3232_),
    .B1(_3081_),
    .B2(_3235_),
    .C1(_3243_),
    .Y(_3244_));
 sky130_fd_sc_hd__and2_1 _3711_ (.A(_3144_),
    .B(_3214_),
    .X(_3245_));
 sky130_fd_sc_hd__clkbuf_2 _3712_ (.A(_3245_),
    .X(_3246_));
 sky130_fd_sc_hd__buf_2 _3713_ (.A(_3246_),
    .X(_3247_));
 sky130_fd_sc_hd__and2_1 _3714_ (.A(_3149_),
    .B(_3215_),
    .X(_3248_));
 sky130_fd_sc_hd__clkbuf_2 _3715_ (.A(_3248_),
    .X(_3249_));
 sky130_fd_sc_hd__clkbuf_4 _3716_ (.A(_3249_),
    .X(_3250_));
 sky130_fd_sc_hd__inv_2 _3717_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_3251_));
 sky130_fd_sc_hd__nand2_2 _3718_ (.A(_3154_),
    .B(_3215_),
    .Y(_3252_));
 sky130_fd_sc_hd__clkbuf_4 _3719_ (.A(_3252_),
    .X(_3253_));
 sky130_fd_sc_hd__and2_1 _3720_ (.A(_3157_),
    .B(_3214_),
    .X(_3254_));
 sky130_fd_sc_hd__clkbuf_2 _3721_ (.A(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__buf_2 _3722_ (.A(_3255_),
    .X(_3256_));
 sky130_fd_sc_hd__nand2_1 _3723_ (.A(_3256_),
    .B(_3056_),
    .Y(_3257_));
 sky130_fd_sc_hd__o21ai_1 _3724_ (.A1(_3251_),
    .A2(_3253_),
    .B1(_3257_),
    .Y(_3258_));
 sky130_fd_sc_hd__a221oi_1 _3725_ (.A1(_3059_),
    .A2(_3247_),
    .B1(_3062_),
    .B2(_3250_),
    .C1(_3258_),
    .Y(_3259_));
 sky130_fd_sc_hd__and2_1 _3726_ (.A(_3191_),
    .B(_3214_),
    .X(_3260_));
 sky130_fd_sc_hd__clkbuf_2 _3727_ (.A(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__clkbuf_4 _3728_ (.A(_3261_),
    .X(_3262_));
 sky130_fd_sc_hd__and2_1 _3729_ (.A(_3010_),
    .B(_3214_),
    .X(_3263_));
 sky130_fd_sc_hd__clkbuf_2 _3730_ (.A(_3263_),
    .X(_3264_));
 sky130_fd_sc_hd__clkbuf_4 _3731_ (.A(_3264_),
    .X(_3265_));
 sky130_fd_sc_hd__inv_2 _3732_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_3266_));
 sky130_fd_sc_hd__nand2_2 _3733_ (.A(_3205_),
    .B(_3215_),
    .Y(_3267_));
 sky130_fd_sc_hd__buf_2 _3734_ (.A(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__inv_2 _3735_ (.A(_3093_),
    .Y(_3269_));
 sky130_fd_sc_hd__nand2_2 _3736_ (.A(_3199_),
    .B(_3215_),
    .Y(_3270_));
 sky130_fd_sc_hd__buf_2 _3737_ (.A(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__o22ai_1 _3738_ (.A1(_3266_),
    .A2(_3268_),
    .B1(_3269_),
    .B2(_3271_),
    .Y(_3272_));
 sky130_fd_sc_hd__a221oi_1 _3739_ (.A1(_3096_),
    .A2(_3262_),
    .B1(_3099_),
    .B2(_3265_),
    .C1(_3272_),
    .Y(_3273_));
 sky130_fd_sc_hd__and4_1 _3740_ (.A(_3229_),
    .B(_3244_),
    .C(_3259_),
    .D(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__buf_2 _3741_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_3275_));
 sky130_fd_sc_hd__or3_2 _3742_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .B(_3011_),
    .C(_3109_),
    .X(_3276_));
 sky130_fd_sc_hd__inv_2 _3743_ (.A(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__clkbuf_4 _3744_ (.A(_3277_),
    .X(_3278_));
 sky130_fd_sc_hd__and2_1 _3745_ (.A(_3108_),
    .B(_3278_),
    .X(_3279_));
 sky130_fd_sc_hd__clkbuf_2 _3746_ (.A(_3279_),
    .X(_3280_));
 sky130_fd_sc_hd__buf_2 _3747_ (.A(_3280_),
    .X(_3281_));
 sky130_fd_sc_hd__buf_2 _3748_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_3282_));
 sky130_fd_sc_hd__and2_1 _3749_ (.A(_3119_),
    .B(_3278_),
    .X(_3283_));
 sky130_fd_sc_hd__clkbuf_2 _3750_ (.A(_3283_),
    .X(_3284_));
 sky130_fd_sc_hd__buf_4 _3751_ (.A(_3284_),
    .X(_3285_));
 sky130_fd_sc_hd__inv_2 _3752_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_3286_));
 sky130_fd_sc_hd__nand2_2 _3753_ (.A(_3128_),
    .B(_3278_),
    .Y(_3287_));
 sky130_fd_sc_hd__buf_2 _3754_ (.A(_3287_),
    .X(_3288_));
 sky130_fd_sc_hd__inv_2 _3755_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_3289_));
 sky130_fd_sc_hd__nand2_2 _3756_ (.A(_3136_),
    .B(_3278_),
    .Y(_3290_));
 sky130_fd_sc_hd__buf_2 _3757_ (.A(_3290_),
    .X(_3291_));
 sky130_fd_sc_hd__o22ai_1 _3758_ (.A1(_3286_),
    .A2(_3288_),
    .B1(_3289_),
    .B2(_3291_),
    .Y(_3292_));
 sky130_fd_sc_hd__a221oi_1 _3759_ (.A1(_3275_),
    .A2(_3281_),
    .B1(_3282_),
    .B2(_3285_),
    .C1(_3292_),
    .Y(_3293_));
 sky130_fd_sc_hd__inv_2 _3760_ (.A(_3157_),
    .Y(_3294_));
 sky130_fd_sc_hd__nor2_2 _3761_ (.A(_3276_),
    .B(_3294_),
    .Y(_3295_));
 sky130_fd_sc_hd__buf_2 _3762_ (.A(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__nand2_1 _3763_ (.A(_3296_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_3297_));
 sky130_fd_sc_hd__and2_1 _3764_ (.A(_3149_),
    .B(_3277_),
    .X(_3298_));
 sky130_fd_sc_hd__clkbuf_2 _3765_ (.A(_3298_),
    .X(_3299_));
 sky130_fd_sc_hd__buf_2 _3766_ (.A(_3299_),
    .X(_3300_));
 sky130_fd_sc_hd__clkbuf_4 _3767_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .X(_3301_));
 sky130_fd_sc_hd__nand2_1 _3768_ (.A(_3300_),
    .B(_3301_),
    .Y(_3302_));
 sky130_fd_sc_hd__and2_1 _3769_ (.A(_3154_),
    .B(_3277_),
    .X(_3303_));
 sky130_fd_sc_hd__clkbuf_2 _3770_ (.A(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__buf_2 _3771_ (.A(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__nand2_1 _3772_ (.A(_3305_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_3306_));
 sky130_fd_sc_hd__and2_1 _3773_ (.A(_3144_),
    .B(_3277_),
    .X(_3307_));
 sky130_fd_sc_hd__clkbuf_2 _3774_ (.A(_3307_),
    .X(_3308_));
 sky130_fd_sc_hd__buf_2 _3775_ (.A(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__nand2_1 _3776_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_3310_));
 sky130_fd_sc_hd__and4_1 _3777_ (.A(_3297_),
    .B(_3302_),
    .C(_3306_),
    .D(_3310_),
    .X(_3311_));
 sky130_fd_sc_hd__inv_2 _3778_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_3312_));
 sky130_fd_sc_hd__nand2_2 _3779_ (.A(_3171_),
    .B(_3278_),
    .Y(_3313_));
 sky130_fd_sc_hd__clkbuf_4 _3780_ (.A(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__inv_2 _3781_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_3315_));
 sky130_fd_sc_hd__nand2_2 _3782_ (.A(_3185_),
    .B(_3278_),
    .Y(_3316_));
 sky130_fd_sc_hd__clkbuf_4 _3783_ (.A(_3316_),
    .X(_3317_));
 sky130_fd_sc_hd__o22ai_1 _3784_ (.A1(_3312_),
    .A2(_3314_),
    .B1(_3315_),
    .B2(_3317_),
    .Y(_3318_));
 sky130_fd_sc_hd__and2_2 _3785_ (.A(_3177_),
    .B(_3278_),
    .X(_3319_));
 sky130_fd_sc_hd__buf_2 _3786_ (.A(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__and2_2 _3787_ (.A(_3167_),
    .B(_3278_),
    .X(_3321_));
 sky130_fd_sc_hd__clkbuf_4 _3788_ (.A(_3321_),
    .X(_3322_));
 sky130_fd_sc_hd__clkbuf_4 _3789_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_3323_));
 sky130_fd_sc_hd__a22o_1 _3790_ (.A1(_3320_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .B1(_3322_),
    .B2(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__nor2_1 _3791_ (.A(_3318_),
    .B(_3324_),
    .Y(_3325_));
 sky130_fd_sc_hd__buf_2 _3792_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .X(_3326_));
 sky130_fd_sc_hd__and2_1 _3793_ (.A(_3191_),
    .B(_3277_),
    .X(_3327_));
 sky130_fd_sc_hd__clkbuf_2 _3794_ (.A(_3327_),
    .X(_3328_));
 sky130_fd_sc_hd__buf_2 _3795_ (.A(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__buf_2 _3796_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .X(_3330_));
 sky130_fd_sc_hd__and2_1 _3797_ (.A(_3010_),
    .B(_3277_),
    .X(_3331_));
 sky130_fd_sc_hd__clkbuf_2 _3798_ (.A(_3331_),
    .X(_3332_));
 sky130_fd_sc_hd__buf_2 _3799_ (.A(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__inv_2 _3800_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_3334_));
 sky130_fd_sc_hd__nand2_2 _3801_ (.A(_3205_),
    .B(_3278_),
    .Y(_3335_));
 sky130_fd_sc_hd__buf_2 _3802_ (.A(_3335_),
    .X(_3336_));
 sky130_fd_sc_hd__inv_2 _3803_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_3337_));
 sky130_fd_sc_hd__nand2_2 _3804_ (.A(_3199_),
    .B(_3278_),
    .Y(_3338_));
 sky130_fd_sc_hd__buf_2 _3805_ (.A(_3338_),
    .X(_3339_));
 sky130_fd_sc_hd__o22ai_1 _3806_ (.A1(_3334_),
    .A2(_3336_),
    .B1(_3337_),
    .B2(_3339_),
    .Y(_3340_));
 sky130_fd_sc_hd__a221oi_1 _3807_ (.A1(_3326_),
    .A2(_3329_),
    .B1(_3330_),
    .B2(_3333_),
    .C1(_3340_),
    .Y(_3341_));
 sky130_fd_sc_hd__and4_1 _3808_ (.A(_3293_),
    .B(_3311_),
    .C(_3325_),
    .D(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__clkbuf_4 _3809_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .X(_3343_));
 sky130_fd_sc_hd__or3_1 _3810_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .B(_3011_),
    .C(_3110_),
    .X(_3344_));
 sky130_fd_sc_hd__inv_2 _3811_ (.A(_3344_),
    .Y(_3345_));
 sky130_fd_sc_hd__buf_2 _3812_ (.A(_3345_),
    .X(_3346_));
 sky130_fd_sc_hd__and2_1 _3813_ (.A(_3108_),
    .B(_3346_),
    .X(_3347_));
 sky130_fd_sc_hd__clkbuf_2 _3814_ (.A(_3347_),
    .X(_3348_));
 sky130_fd_sc_hd__buf_2 _3815_ (.A(_3348_),
    .X(_3349_));
 sky130_fd_sc_hd__buf_2 _3816_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .X(_3350_));
 sky130_fd_sc_hd__and2_1 _3817_ (.A(_3119_),
    .B(_3346_),
    .X(_3351_));
 sky130_fd_sc_hd__clkbuf_2 _3818_ (.A(_3351_),
    .X(_3352_));
 sky130_fd_sc_hd__buf_4 _3819_ (.A(_3352_),
    .X(_3353_));
 sky130_fd_sc_hd__and2_1 _3820_ (.A(_3136_),
    .B(_3346_),
    .X(_3354_));
 sky130_fd_sc_hd__clkbuf_2 _3821_ (.A(_3354_),
    .X(_3355_));
 sky130_fd_sc_hd__buf_6 _3822_ (.A(_3355_),
    .X(_3356_));
 sky130_fd_sc_hd__clkbuf_4 _3823_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .X(_3357_));
 sky130_fd_sc_hd__nand2_1 _3824_ (.A(_3356_),
    .B(_3357_),
    .Y(_3358_));
 sky130_fd_sc_hd__and2_1 _3825_ (.A(_3128_),
    .B(_3346_),
    .X(_3359_));
 sky130_fd_sc_hd__clkbuf_2 _3826_ (.A(_3359_),
    .X(_3360_));
 sky130_fd_sc_hd__buf_2 _3827_ (.A(_3360_),
    .X(_3361_));
 sky130_fd_sc_hd__clkbuf_4 _3828_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .X(_3362_));
 sky130_fd_sc_hd__nand2_1 _3829_ (.A(_3361_),
    .B(_3362_),
    .Y(_3363_));
 sky130_fd_sc_hd__nand2_1 _3830_ (.A(_3358_),
    .B(_3363_),
    .Y(_3364_));
 sky130_fd_sc_hd__a221oi_1 _3831_ (.A1(_3343_),
    .A2(_3349_),
    .B1(_3350_),
    .B2(_3353_),
    .C1(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__buf_2 _3832_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .X(_3366_));
 sky130_fd_sc_hd__and2_1 _3833_ (.A(_3154_),
    .B(_3346_),
    .X(_3367_));
 sky130_fd_sc_hd__clkbuf_2 _3834_ (.A(_3367_),
    .X(_3368_));
 sky130_fd_sc_hd__buf_2 _3835_ (.A(_3368_),
    .X(_3369_));
 sky130_fd_sc_hd__clkbuf_4 _3836_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .X(_3370_));
 sky130_fd_sc_hd__nor2_2 _3837_ (.A(_3344_),
    .B(_3294_),
    .Y(_3371_));
 sky130_fd_sc_hd__buf_2 _3838_ (.A(_3371_),
    .X(_3372_));
 sky130_fd_sc_hd__and2_1 _3839_ (.A(_3149_),
    .B(_3345_),
    .X(_3373_));
 sky130_fd_sc_hd__clkbuf_2 _3840_ (.A(_3373_),
    .X(_3374_));
 sky130_fd_sc_hd__buf_2 _3841_ (.A(_3374_),
    .X(_3375_));
 sky130_fd_sc_hd__buf_2 _3842_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .X(_3376_));
 sky130_fd_sc_hd__nand2_1 _3843_ (.A(_3375_),
    .B(_3376_),
    .Y(_3377_));
 sky130_fd_sc_hd__and2_1 _3844_ (.A(_3144_),
    .B(_3345_),
    .X(_3378_));
 sky130_fd_sc_hd__clkbuf_2 _3845_ (.A(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__buf_2 _3846_ (.A(_3379_),
    .X(_3380_));
 sky130_fd_sc_hd__buf_2 _3847_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .X(_3381_));
 sky130_fd_sc_hd__nand2_1 _3848_ (.A(_3380_),
    .B(_3381_),
    .Y(_3382_));
 sky130_fd_sc_hd__nand2_1 _3849_ (.A(_3377_),
    .B(_3382_),
    .Y(_3383_));
 sky130_fd_sc_hd__a221oi_1 _3850_ (.A1(_3366_),
    .A2(_3369_),
    .B1(_3370_),
    .B2(_3372_),
    .C1(_3383_),
    .Y(_3384_));
 sky130_fd_sc_hd__inv_2 _3851_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_3385_));
 sky130_fd_sc_hd__nand2_2 _3852_ (.A(_3167_),
    .B(_3346_),
    .Y(_3386_));
 sky130_fd_sc_hd__buf_2 _3853_ (.A(_3386_),
    .X(_3387_));
 sky130_fd_sc_hd__and2_1 _3854_ (.A(_3171_),
    .B(_3345_),
    .X(_3388_));
 sky130_fd_sc_hd__clkbuf_2 _3855_ (.A(_3388_),
    .X(_3389_));
 sky130_fd_sc_hd__buf_4 _3856_ (.A(_3389_),
    .X(_3390_));
 sky130_fd_sc_hd__clkbuf_4 _3857_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_3391_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_3390_),
    .B(_3391_),
    .Y(_3392_));
 sky130_fd_sc_hd__and2_1 _3859_ (.A(_3177_),
    .B(_3345_),
    .X(_3393_));
 sky130_fd_sc_hd__clkbuf_2 _3860_ (.A(_3393_),
    .X(_3394_));
 sky130_fd_sc_hd__buf_2 _3861_ (.A(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__buf_2 _3862_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .X(_3396_));
 sky130_fd_sc_hd__nand2_1 _3863_ (.A(_3395_),
    .B(_3396_),
    .Y(_3397_));
 sky130_fd_sc_hd__inv_2 _3864_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_3398_));
 sky130_fd_sc_hd__nand2_2 _3865_ (.A(_3185_),
    .B(_3346_),
    .Y(_3399_));
 sky130_fd_sc_hd__clkbuf_2 _3866_ (.A(_3399_),
    .X(_3400_));
 sky130_fd_sc_hd__or2_1 _3867_ (.A(_3398_),
    .B(_3400_),
    .X(_3401_));
 sky130_fd_sc_hd__o2111a_1 _3868_ (.A1(_3385_),
    .A2(_3387_),
    .B1(_3392_),
    .C1(_3397_),
    .D1(_3401_),
    .X(_3402_));
 sky130_fd_sc_hd__buf_2 _3869_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .X(_3403_));
 sky130_fd_sc_hd__and2_1 _3870_ (.A(_3205_),
    .B(_3346_),
    .X(_3404_));
 sky130_fd_sc_hd__clkbuf_2 _3871_ (.A(_3404_),
    .X(_3405_));
 sky130_fd_sc_hd__clkbuf_4 _3872_ (.A(_3405_),
    .X(_3406_));
 sky130_fd_sc_hd__buf_2 _3873_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .X(_3407_));
 sky130_fd_sc_hd__and2_1 _3874_ (.A(_3199_),
    .B(_3346_),
    .X(_3408_));
 sky130_fd_sc_hd__clkbuf_2 _3875_ (.A(_3408_),
    .X(_3409_));
 sky130_fd_sc_hd__clkbuf_4 _3876_ (.A(_3409_),
    .X(_3410_));
 sky130_fd_sc_hd__inv_2 _3877_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_3411_));
 sky130_fd_sc_hd__nand2_2 _3878_ (.A(_3010_),
    .B(_3346_),
    .Y(_3412_));
 sky130_fd_sc_hd__clkbuf_4 _3879_ (.A(_3412_),
    .X(_3413_));
 sky130_fd_sc_hd__and2_1 _3880_ (.A(_3191_),
    .B(_3345_),
    .X(_3414_));
 sky130_fd_sc_hd__clkbuf_2 _3881_ (.A(_3414_),
    .X(_3415_));
 sky130_fd_sc_hd__buf_2 _3882_ (.A(_3415_),
    .X(_3416_));
 sky130_fd_sc_hd__nand2_1 _3883_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_3417_));
 sky130_fd_sc_hd__o21ai_1 _3884_ (.A1(_3411_),
    .A2(_3413_),
    .B1(_3417_),
    .Y(_0322_));
 sky130_fd_sc_hd__a221oi_1 _3885_ (.A1(_3403_),
    .A2(_3406_),
    .B1(_3407_),
    .B2(_3410_),
    .C1(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__and4_1 _3886_ (.A(_3365_),
    .B(_3384_),
    .C(_3402_),
    .D(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__and4_1 _3887_ (.A(_3213_),
    .B(_3274_),
    .C(_3342_),
    .D(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_4 _3888_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_0326_));
 sky130_fd_sc_hd__and3_2 _3889_ (.A(_3011_),
    .B(_3109_),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_0327_));
 sky130_fd_sc_hd__buf_2 _3890_ (.A(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__and2_1 _3891_ (.A(_3108_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_2 _3892_ (.A(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__buf_2 _3893_ (.A(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__buf_2 _3894_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_0332_));
 sky130_fd_sc_hd__and2_1 _3895_ (.A(_3119_),
    .B(_0328_),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_2 _3896_ (.A(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__buf_6 _3897_ (.A(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__and2_1 _3898_ (.A(_3136_),
    .B(_0327_),
    .X(_0336_));
 sky130_fd_sc_hd__buf_6 _3899_ (.A(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__buf_6 _3900_ (.A(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_4 _3901_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _3902_ (.A(_0338_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__and2_1 _3903_ (.A(_3128_),
    .B(_0327_),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_2 _3904_ (.A(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__buf_4 _3905_ (.A(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_4 _3906_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_0344_));
 sky130_fd_sc_hd__nand2_1 _3907_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_0340_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a221oi_1 _3909_ (.A1(_0326_),
    .A2(_0331_),
    .B1(_0332_),
    .B2(_0335_),
    .C1(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _3910_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_2 _3911_ (.A(_3171_),
    .B(_0328_),
    .Y(_0349_));
 sky130_fd_sc_hd__clkbuf_4 _3912_ (.A(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__inv_2 _3913_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_2 _3914_ (.A(_3185_),
    .B(_0328_),
    .Y(_0352_));
 sky130_fd_sc_hd__buf_2 _3915_ (.A(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__o22ai_1 _3916_ (.A1(_0348_),
    .A2(_0350_),
    .B1(_0351_),
    .B2(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__and2_2 _3917_ (.A(_3177_),
    .B(_0328_),
    .X(_0355_));
 sky130_fd_sc_hd__buf_2 _3918_ (.A(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_4 _3919_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_0357_));
 sky130_fd_sc_hd__and2_2 _3920_ (.A(_3167_),
    .B(_0328_),
    .X(_0358_));
 sky130_fd_sc_hd__buf_2 _3921_ (.A(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__buf_2 _3922_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _3923_ (.A1(_0356_),
    .A2(_0357_),
    .B1(_0359_),
    .B2(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__nor2_1 _3924_ (.A(_0354_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__clkbuf_4 _3925_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _3926_ (.A(_3154_),
    .B(_0327_),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_2 _3927_ (.A(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_2 _3928_ (.A(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__buf_2 _3929_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _3930_ (.A(_3157_),
    .B(_0328_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_2 _3931_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__buf_2 _3932_ (.A(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__inv_2 _3933_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_2 _3934_ (.A(_3144_),
    .B(_0328_),
    .Y(_0372_));
 sky130_fd_sc_hd__clkbuf_4 _3935_ (.A(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__and2_1 _3936_ (.A(_3149_),
    .B(_0327_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_2 _3937_ (.A(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__buf_2 _3938_ (.A(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_4 _3939_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _3940_ (.A(_0376_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__o21ai_1 _3941_ (.A1(_0371_),
    .A2(_0373_),
    .B1(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__a221oi_1 _3942_ (.A1(_0363_),
    .A2(_0366_),
    .B1(_0367_),
    .B2(_0370_),
    .C1(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__buf_2 _3943_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _3944_ (.A(_3205_),
    .B(_0327_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_2 _3945_ (.A(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_4 _3946_ (.A(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__buf_2 _3947_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _3948_ (.A(_3199_),
    .B(_0328_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_2 _3949_ (.A(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_2 _3950_ (.A(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__inv_2 _3951_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_2 _3952_ (.A(_3010_),
    .B(_0328_),
    .Y(_0390_));
 sky130_fd_sc_hd__clkbuf_4 _3953_ (.A(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__and2_1 _3954_ (.A(_3191_),
    .B(_0327_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_2 _3955_ (.A(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__buf_2 _3956_ (.A(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _3957_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_0395_));
 sky130_fd_sc_hd__o21ai_1 _3958_ (.A1(_0389_),
    .A2(_0391_),
    .B1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__a221oi_1 _3959_ (.A1(_0381_),
    .A2(_0384_),
    .B1(_0385_),
    .B2(_0388_),
    .C1(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__and4_1 _3960_ (.A(_0347_),
    .B(_0362_),
    .C(_0380_),
    .D(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__inv_2 _3961_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_0399_));
 sky130_fd_sc_hd__buf_2 _3962_ (.A(_3012_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_2 _3963_ (.A(_3185_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__buf_2 _3964_ (.A(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__and2_1 _3965_ (.A(_3177_),
    .B(_3012_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_2 _3966_ (.A(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__buf_2 _3967_ (.A(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_1 _3968_ (.A(_0405_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0406_));
 sky130_fd_sc_hd__and2_1 _3969_ (.A(_3171_),
    .B(_0400_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_2 _3970_ (.A(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__buf_4 _3971_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__buf_2 _3972_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_0410_));
 sky130_fd_sc_hd__nand2_1 _3973_ (.A(_0409_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__inv_2 _3974_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _3975_ (.A(_3167_),
    .B(_0400_),
    .Y(_0413_));
 sky130_fd_sc_hd__clkbuf_2 _3976_ (.A(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__or2_1 _3977_ (.A(_0412_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__o2111a_1 _3978_ (.A1(_0399_),
    .A2(_0402_),
    .B1(_0406_),
    .C1(_0411_),
    .D1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__inv_2 _3979_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .Y(_0417_));
 sky130_fd_sc_hd__nand2_2 _3980_ (.A(_3119_),
    .B(_0400_),
    .Y(_0418_));
 sky130_fd_sc_hd__buf_2 _3981_ (.A(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__and2_1 _3982_ (.A(_3128_),
    .B(_3012_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_2 _3983_ (.A(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__buf_4 _3984_ (.A(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _3985_ (.A(_0422_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0423_));
 sky130_fd_sc_hd__and2_1 _3986_ (.A(_3108_),
    .B(_3012_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_2 _3987_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__buf_2 _3988_ (.A(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__buf_2 _3989_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _3990_ (.A(_0426_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _3991_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0429_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(_3136_),
    .B(_0400_),
    .Y(_0430_));
 sky130_fd_sc_hd__buf_2 _3993_ (.A(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__or2_1 _3994_ (.A(_0429_),
    .B(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__o2111a_1 _3995_ (.A1(_0417_),
    .A2(_0419_),
    .B1(_0423_),
    .C1(_0428_),
    .D1(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__buf_2 _3996_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_0434_));
 sky130_fd_sc_hd__and2_1 _3997_ (.A(_3144_),
    .B(_0400_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_2 _3998_ (.A(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__buf_2 _3999_ (.A(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__buf_2 _4000_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_0438_));
 sky130_fd_sc_hd__and2_1 _4001_ (.A(_3149_),
    .B(_0400_),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_2 _4002_ (.A(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__buf_2 _4003_ (.A(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__inv_2 _4004_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_2 _4005_ (.A(_3154_),
    .B(_0400_),
    .Y(_0443_));
 sky130_fd_sc_hd__clkbuf_4 _4006_ (.A(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__and2_1 _4007_ (.A(_3157_),
    .B(_3012_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_2 _4008_ (.A(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__buf_2 _4009_ (.A(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__buf_2 _4010_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_0448_));
 sky130_fd_sc_hd__nand2_1 _4011_ (.A(_0447_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__o21ai_1 _4012_ (.A1(_0442_),
    .A2(_0444_),
    .B1(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__a221oi_1 _4013_ (.A1(_0434_),
    .A2(_0437_),
    .B1(_0438_),
    .B2(_0441_),
    .C1(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _4014_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .X(_0452_));
 sky130_fd_sc_hd__and2_1 _4015_ (.A(_3205_),
    .B(_0400_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_2 _4016_ (.A(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__buf_2 _4017_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__buf_2 _4018_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .X(_0456_));
 sky130_fd_sc_hd__and2_1 _4019_ (.A(_3199_),
    .B(_0400_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_2 _4020_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_4 _4021_ (.A(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__inv_2 _4022_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_0460_));
 sky130_fd_sc_hd__inv_2 _4023_ (.A(_3013_),
    .Y(_0461_));
 sky130_fd_sc_hd__clkbuf_4 _4024_ (.A(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__and2_1 _4025_ (.A(_3191_),
    .B(_3012_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_2 _4026_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__buf_2 _4027_ (.A(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__nand2_1 _4028_ (.A(_0465_),
    .B(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_0466_));
 sky130_fd_sc_hd__o21ai_1 _4029_ (.A1(_0460_),
    .A2(_0462_),
    .B1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__a221oi_1 _4030_ (.A1(_0452_),
    .A2(_0455_),
    .B1(_0456_),
    .B2(_0459_),
    .C1(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__and4_1 _4031_ (.A(_0416_),
    .B(_0433_),
    .C(_0451_),
    .D(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__and2_1 _4032_ (.A(_0398_),
    .B(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_4 _4033_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .X(_0471_));
 sky130_fd_sc_hd__inv_2 _4034_ (.A(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__and3_2 _4035_ (.A(_3011_),
    .B(_3110_),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_0473_));
 sky130_fd_sc_hd__buf_2 _4036_ (.A(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__nand2_2 _4037_ (.A(_3128_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__buf_2 _4038_ (.A(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__and2_1 _4039_ (.A(_3136_),
    .B(_0474_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_2 _4040_ (.A(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_2 _4041_ (.A(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_4 _4042_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .X(_0480_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(_0479_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__and2_2 _4044_ (.A(_3108_),
    .B(_0473_),
    .X(_0482_));
 sky130_fd_sc_hd__buf_2 _4045_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__and2_2 _4046_ (.A(_3119_),
    .B(_0473_),
    .X(_0484_));
 sky130_fd_sc_hd__buf_2 _4047_ (.A(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_4 _4048_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_1 _4049_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .B1(_0485_),
    .B2(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__inv_2 _4050_ (.A(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__o211a_1 _4051_ (.A1(_0472_),
    .A2(_0476_),
    .B1(_0481_),
    .C1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__and2_1 _4052_ (.A(_3154_),
    .B(_0474_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_2 _4053_ (.A(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__buf_2 _4054_ (.A(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_4 _4055_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _4056_ (.A(_3157_),
    .B(_0474_),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_2 _4057_ (.A(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__buf_2 _4058_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_4 _4059_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .X(_0497_));
 sky130_fd_sc_hd__inv_2 _4060_ (.A(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2_2 _4061_ (.A(_3144_),
    .B(_0474_),
    .Y(_0499_));
 sky130_fd_sc_hd__clkbuf_4 _4062_ (.A(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__and2_1 _4063_ (.A(_3149_),
    .B(_0474_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_2 _4064_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__buf_2 _4065_ (.A(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_4 _4066_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_1 _4067_ (.A(_0503_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__o21ai_1 _4068_ (.A1(_0498_),
    .A2(_0500_),
    .B1(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__a221oi_1 _4069_ (.A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .A2(_0492_),
    .B1(_0493_),
    .B2(_0496_),
    .C1(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__clkbuf_4 _4070_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .X(_0508_));
 sky130_fd_sc_hd__inv_2 _4071_ (.A(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_2 _4072_ (.A(_3167_),
    .B(_0474_),
    .Y(_0510_));
 sky130_fd_sc_hd__buf_2 _4073_ (.A(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__and2_1 _4074_ (.A(_3177_),
    .B(_0473_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_2 _4075_ (.A(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__buf_2 _4076_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _4077_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _4078_ (.A(_0514_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__and2_1 _4079_ (.A(_3171_),
    .B(_0473_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_2 _4080_ (.A(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__buf_2 _4081_ (.A(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_4 _4082_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(_0519_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__clkbuf_4 _4084_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .X(_0522_));
 sky130_fd_sc_hd__inv_2 _4085_ (.A(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2_2 _4086_ (.A(_3185_),
    .B(_0474_),
    .Y(_0524_));
 sky130_fd_sc_hd__clkbuf_2 _4087_ (.A(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_1 _4088_ (.A(_0523_),
    .B(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__o2111a_1 _4089_ (.A1(_0509_),
    .A2(_0511_),
    .B1(_0516_),
    .C1(_0521_),
    .D1(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _4090_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_0528_));
 sky130_fd_sc_hd__and2_1 _4091_ (.A(_3191_),
    .B(_0474_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_2 _4092_ (.A(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__buf_2 _4093_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_4 _4094_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_0532_));
 sky130_fd_sc_hd__and2_1 _4095_ (.A(_3010_),
    .B(_0474_),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_2 _4096_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__buf_2 _4097_ (.A(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__and2_1 _4098_ (.A(_3199_),
    .B(_0473_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_2 _4099_ (.A(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_2 _4100_ (.A(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__buf_2 _4101_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_1 _4102_ (.A(_0538_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__and2_1 _4103_ (.A(_3205_),
    .B(_0473_),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_2 _4104_ (.A(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__buf_2 _4105_ (.A(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_4 _4106_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_1 _4107_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _4108_ (.A(_0540_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__a221oi_1 _4109_ (.A1(_0528_),
    .A2(_0531_),
    .B1(_0532_),
    .B2(_0535_),
    .C1(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__and4_1 _4110_ (.A(_0489_),
    .B(_0507_),
    .C(_0527_),
    .D(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_4 _4111_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_0549_));
 sky130_fd_sc_hd__inv_2 _4112_ (.A(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__and3_2 _4113_ (.A(_3011_),
    .B(_3109_),
    .C(_3110_),
    .X(_0551_));
 sky130_fd_sc_hd__buf_4 _4114_ (.A(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_2 _4115_ (.A(_3185_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__clkbuf_4 _4116_ (.A(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__and2_1 _4117_ (.A(_3177_),
    .B(_0551_),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_2 _4118_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__buf_2 _4119_ (.A(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_4 _4120_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _4121_ (.A(_0557_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__and2_1 _4122_ (.A(_3171_),
    .B(_0551_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_2 _4123_ (.A(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__buf_2 _4124_ (.A(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_4 _4125_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_1 _4126_ (.A(_0562_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__inv_2 _4127_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_2 _4128_ (.A(_3167_),
    .B(_0552_),
    .Y(_0566_));
 sky130_fd_sc_hd__clkbuf_2 _4129_ (.A(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__or2_1 _4130_ (.A(_0565_),
    .B(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__o2111a_1 _4131_ (.A1(_0550_),
    .A2(_0554_),
    .B1(_0559_),
    .C1(_0564_),
    .D1(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__inv_2 _4132_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_2 _4133_ (.A(_3119_),
    .B(_0552_),
    .Y(_0571_));
 sky130_fd_sc_hd__buf_2 _4134_ (.A(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__and2_1 _4135_ (.A(_3108_),
    .B(_0551_),
    .X(_0573_));
 sky130_fd_sc_hd__clkbuf_2 _4136_ (.A(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__buf_2 _4137_ (.A(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_1 _4138_ (.A(_0575_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0576_));
 sky130_fd_sc_hd__and2_1 _4139_ (.A(_3128_),
    .B(_0551_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_2 _4140_ (.A(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__buf_2 _4141_ (.A(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__nand2_1 _4142_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_2 _4143_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_2 _4144_ (.A(_3136_),
    .B(_0552_),
    .Y(_0582_));
 sky130_fd_sc_hd__clkbuf_2 _4145_ (.A(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__or2_1 _4146_ (.A(_0581_),
    .B(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__o2111a_1 _4147_ (.A1(_0570_),
    .A2(_0572_),
    .B1(_0576_),
    .C1(_0580_),
    .D1(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_4 _4148_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_0586_));
 sky130_fd_sc_hd__inv_2 _4149_ (.A(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__nand2_2 _4150_ (.A(_3144_),
    .B(_0552_),
    .Y(_0588_));
 sky130_fd_sc_hd__buf_2 _4151_ (.A(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__inv_2 _4152_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_2 _4153_ (.A(_3157_),
    .B(_0552_),
    .Y(_0591_));
 sky130_fd_sc_hd__buf_2 _4154_ (.A(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_4 _4155_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_0593_));
 sky130_fd_sc_hd__inv_2 _4156_ (.A(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _4157_ (.A(_3149_),
    .B(_0552_),
    .Y(_0595_));
 sky130_fd_sc_hd__clkbuf_2 _4158_ (.A(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__or2_1 _4159_ (.A(_0594_),
    .B(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__o221a_1 _4160_ (.A1(_0587_),
    .A2(_0589_),
    .B1(_0590_),
    .B2(_0592_),
    .C1(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__and2_1 _4161_ (.A(_3191_),
    .B(_0551_),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_2 _4162_ (.A(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__buf_2 _4163_ (.A(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__and2_1 _4164_ (.A(_3010_),
    .B(_0551_),
    .X(_0602_));
 sky130_fd_sc_hd__clkbuf_2 _4165_ (.A(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__buf_2 _4166_ (.A(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__inv_2 _4167_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_2 _4168_ (.A(_3205_),
    .B(_0552_),
    .Y(_0606_));
 sky130_fd_sc_hd__buf_2 _4169_ (.A(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__inv_2 _4170_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_2 _4171_ (.A(_3199_),
    .B(_0552_),
    .Y(_0609_));
 sky130_fd_sc_hd__buf_2 _4172_ (.A(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__o22ai_1 _4173_ (.A1(_0605_),
    .A2(_0607_),
    .B1(_0608_),
    .B2(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__a221oi_1 _4174_ (.A1(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .A2(_0601_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .B2(_0604_),
    .C1(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__and4_1 _4175_ (.A(_0569_),
    .B(_0585_),
    .C(_0598_),
    .D(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _4176_ (.A(_0470_),
    .B(_0548_),
    .C(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__o41a_1 _4177_ (.A1(\egd_top.BitStream_buffer.pc[2] ),
    .A2(\egd_top.BitStream_buffer.pc[3] ),
    .A3(\egd_top.BitStream_buffer.pc[1] ),
    .A4(_3008_),
    .B1(_0552_),
    .X(_0615_));
 sky130_fd_sc_hd__and4b_1 _4178_ (.A_N(_0615_),
    .B(_3011_),
    .C(_3109_),
    .D(_3110_),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_2 _4179_ (.A(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__clkbuf_4 _4180_ (.A(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__buf_2 _4181_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0619_));
 sky130_fd_sc_hd__nand2_1 _4182_ (.A(_0618_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nand3_1 _4183_ (.A(_0325_),
    .B(_0614_),
    .C(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__o21a_1 _4184_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .A2(_3043_),
    .B1(_2980_),
    .X(_0622_));
 sky130_fd_sc_hd__o21a_1 _4185_ (.A1(_3103_),
    .A2(_0621_),
    .B1(_0622_),
    .X(_0297_));
 sky130_fd_sc_hd__inv_2 _4186_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_0623_));
 sky130_fd_sc_hd__o22ai_1 _4187_ (.A1(_3132_),
    .A2(_3130_),
    .B1(_0623_),
    .B2(_3138_),
    .Y(_0624_));
 sky130_fd_sc_hd__a221oi_1 _4188_ (.A1(_3116_),
    .A2(_3115_),
    .B1(_3209_),
    .B2(_3122_),
    .C1(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_2 _4189_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _4190_ (.A(_3160_),
    .B(_3141_),
    .Y(_0627_));
 sky130_fd_sc_hd__o21ai_1 _4191_ (.A1(_0626_),
    .A2(_3156_),
    .B1(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__a221oi_1 _4192_ (.A1(_3148_),
    .A2(_3147_),
    .B1(_3175_),
    .B2(_3152_),
    .C1(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__buf_2 _4193_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_0630_));
 sky130_fd_sc_hd__nand2_1 _4194_ (.A(_3174_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__buf_2 _4195_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_0632_));
 sky130_fd_sc_hd__nand2_1 _4196_ (.A(_3180_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_0634_));
 sky130_fd_sc_hd__or2_1 _4198_ (.A(_0634_),
    .B(_3187_),
    .X(_0635_));
 sky130_fd_sc_hd__o2111a_1 _4199_ (.A1(_3123_),
    .A2(_3169_),
    .B1(_0631_),
    .C1(_0633_),
    .D1(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_4 _4200_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_0637_));
 sky130_fd_sc_hd__nand2_1 _4201_ (.A(_3202_),
    .B(_3190_),
    .Y(_0638_));
 sky130_fd_sc_hd__nand2_1 _4202_ (.A(_3208_),
    .B(_3203_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _4203_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__a221oi_1 _4204_ (.A1(_3195_),
    .A2(_3194_),
    .B1(_0637_),
    .B2(_3198_),
    .C1(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__and4_1 _4205_ (.A(_0625_),
    .B(_0629_),
    .C(_0636_),
    .D(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__inv_2 _4206_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_0643_));
 sky130_fd_sc_hd__o22ai_1 _4207_ (.A1(_3225_),
    .A2(_3224_),
    .B1(_0643_),
    .B2(_3227_),
    .Y(_0644_));
 sky130_fd_sc_hd__a221oi_1 _4208_ (.A1(_3074_),
    .A2(_3218_),
    .B1(_3078_),
    .B2(_3221_),
    .C1(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _4209_ (.A(_3241_),
    .B(_3087_),
    .Y(_0646_));
 sky130_fd_sc_hd__o21ai_1 _4210_ (.A1(_3266_),
    .A2(_3238_),
    .B1(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__a221oi_1 _4211_ (.A1(_3081_),
    .A2(_3232_),
    .B1(_3084_),
    .B2(_3235_),
    .C1(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__inv_2 _4212_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _4213_ (.A(_3256_),
    .B(_3059_),
    .Y(_0650_));
 sky130_fd_sc_hd__o21ai_1 _4214_ (.A1(_0649_),
    .A2(_3253_),
    .B1(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__a221oi_1 _4215_ (.A1(_3062_),
    .A2(_3247_),
    .B1(_3065_),
    .B2(_3250_),
    .C1(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _4216_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_0653_));
 sky130_fd_sc_hd__o22ai_1 _4217_ (.A1(_3269_),
    .A2(_3268_),
    .B1(_0653_),
    .B2(_3271_),
    .Y(_0654_));
 sky130_fd_sc_hd__a221oi_1 _4218_ (.A1(_3099_),
    .A2(_3262_),
    .B1(_0619_),
    .B2(_3265_),
    .C1(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__and4_1 _4219_ (.A(_0645_),
    .B(_0648_),
    .C(_0652_),
    .D(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_4 _4220_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_0657_));
 sky130_fd_sc_hd__inv_2 _4221_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_0658_));
 sky130_fd_sc_hd__o22ai_1 _4222_ (.A1(_3289_),
    .A2(_3288_),
    .B1(_0658_),
    .B2(_3291_),
    .Y(_0659_));
 sky130_fd_sc_hd__a221oi_1 _4223_ (.A1(_3282_),
    .A2(_3281_),
    .B1(_0657_),
    .B2(_3285_),
    .C1(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__clkbuf_4 _4224_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .X(_0661_));
 sky130_fd_sc_hd__nand2_1 _4225_ (.A(_3296_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__clkbuf_4 _4226_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .X(_0663_));
 sky130_fd_sc_hd__nand2_1 _4227_ (.A(_3300_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(_3305_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _4229_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0666_));
 sky130_fd_sc_hd__and4_1 _4230_ (.A(_0662_),
    .B(_0664_),
    .C(_0665_),
    .D(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__inv_2 _4231_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0668_));
 sky130_fd_sc_hd__o22ai_1 _4232_ (.A1(_3315_),
    .A2(_3314_),
    .B1(_0668_),
    .B2(_3317_),
    .Y(_0669_));
 sky130_fd_sc_hd__clkbuf_4 _4233_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_0670_));
 sky130_fd_sc_hd__a22o_1 _4234_ (.A1(_3320_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .B1(_3322_),
    .B2(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__nor2_1 _4235_ (.A(_0669_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__inv_2 _4236_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_0673_));
 sky130_fd_sc_hd__o22ai_1 _4237_ (.A1(_3337_),
    .A2(_3336_),
    .B1(_0673_),
    .B2(_3339_),
    .Y(_0674_));
 sky130_fd_sc_hd__a221oi_1 _4238_ (.A1(_3330_),
    .A2(_3329_),
    .B1(_3366_),
    .B2(_3333_),
    .C1(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__and4_1 _4239_ (.A(_0660_),
    .B(_0667_),
    .C(_0672_),
    .D(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _4240_ (.A(_3356_),
    .B(_3343_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(_3361_),
    .B(_3357_),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _4242_ (.A(_0677_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__a221oi_1 _4243_ (.A1(_3350_),
    .A2(_3349_),
    .B1(_3403_),
    .B2(_3353_),
    .C1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _4244_ (.A(_3375_),
    .B(_3391_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _4245_ (.A(_3380_),
    .B(_3376_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _4246_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a221oi_1 _4247_ (.A1(_3370_),
    .A2(_3369_),
    .B1(_3381_),
    .B2(_3372_),
    .C1(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _4248_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0685_));
 sky130_fd_sc_hd__buf_2 _4249_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_0686_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(_3390_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__buf_2 _4251_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_1 _4252_ (.A(_3395_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__inv_2 _4253_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_0690_));
 sky130_fd_sc_hd__or2_1 _4254_ (.A(_0690_),
    .B(_3400_),
    .X(_0691_));
 sky130_fd_sc_hd__o2111a_1 _4255_ (.A1(_0685_),
    .A2(_3387_),
    .B1(_0687_),
    .C1(_0689_),
    .D1(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_4 _4256_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .X(_0693_));
 sky130_fd_sc_hd__nand2_1 _4257_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_0694_));
 sky130_fd_sc_hd__o21ai_1 _4258_ (.A1(_3251_),
    .A2(_3413_),
    .B1(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__a221oi_1 _4259_ (.A1(_3407_),
    .A2(_3406_),
    .B1(_0693_),
    .B2(_3410_),
    .C1(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__and4_1 _4260_ (.A(_0680_),
    .B(_0684_),
    .C(_0692_),
    .D(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__and4_1 _4261_ (.A(_0642_),
    .B(_0656_),
    .C(_0676_),
    .D(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__nand2_1 _4262_ (.A(_0338_),
    .B(_0326_),
    .Y(_0699_));
 sky130_fd_sc_hd__nand2_1 _4263_ (.A(_0343_),
    .B(_0339_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand2_1 _4264_ (.A(_0699_),
    .B(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__a221oi_1 _4265_ (.A1(_0332_),
    .A2(_0331_),
    .B1(_0381_),
    .B2(_0335_),
    .C1(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__inv_2 _4266_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .Y(_0703_));
 sky130_fd_sc_hd__o22ai_1 _4267_ (.A1(_0351_),
    .A2(_0350_),
    .B1(_0703_),
    .B2(_0353_),
    .Y(_0704_));
 sky130_fd_sc_hd__a22o_1 _4268_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .B1(_0359_),
    .B2(_0344_),
    .X(_0705_));
 sky130_fd_sc_hd__nor2_1 _4269_ (.A(_0704_),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__buf_2 _4270_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_0707_));
 sky130_fd_sc_hd__inv_2 _4271_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_0708_));
 sky130_fd_sc_hd__clkbuf_4 _4272_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_0709_));
 sky130_fd_sc_hd__nand2_1 _4273_ (.A(_0376_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o21ai_1 _4274_ (.A1(_0708_),
    .A2(_0373_),
    .B1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__a221oi_1 _4275_ (.A1(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .A2(_0366_),
    .B1(_0707_),
    .B2(_0370_),
    .C1(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__buf_2 _4276_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_0713_));
 sky130_fd_sc_hd__buf_2 _4277_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_1 _4278_ (.A(_0394_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__o21ai_1 _4279_ (.A1(_0442_),
    .A2(_0391_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a221oi_1 _4280_ (.A1(_0385_),
    .A2(_0384_),
    .B1(_0713_),
    .B2(_0388_),
    .C1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__and4_1 _4281_ (.A(_0702_),
    .B(_0706_),
    .C(_0712_),
    .D(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__inv_2 _4282_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0719_));
 sky130_fd_sc_hd__buf_2 _4283_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .X(_0720_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_0405_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__buf_2 _4285_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(_0409_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__inv_2 _4287_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0724_));
 sky130_fd_sc_hd__or2_1 _4288_ (.A(_0724_),
    .B(_0414_),
    .X(_0725_));
 sky130_fd_sc_hd__o2111a_1 _4289_ (.A1(_0719_),
    .A2(_0402_),
    .B1(_0721_),
    .C1(_0723_),
    .D1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__inv_2 _4290_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _4291_ (.A(_0422_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0728_));
 sky130_fd_sc_hd__buf_2 _4292_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .X(_0729_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(_0426_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__inv_2 _4294_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0731_));
 sky130_fd_sc_hd__or2_1 _4295_ (.A(_0731_),
    .B(_0431_),
    .X(_0732_));
 sky130_fd_sc_hd__o2111a_1 _4296_ (.A1(_0727_),
    .A2(_0419_),
    .B1(_0728_),
    .C1(_0730_),
    .D1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__inv_2 _4297_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_0447_),
    .B(_0434_),
    .Y(_0735_));
 sky130_fd_sc_hd__o21ai_1 _4299_ (.A1(_0734_),
    .A2(_0444_),
    .B1(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__a221oi_1 _4300_ (.A1(_0438_),
    .A2(_0437_),
    .B1(_0410_),
    .B2(_0441_),
    .C1(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__buf_2 _4301_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .X(_0738_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_0465_),
    .B(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_0739_));
 sky130_fd_sc_hd__o21ai_1 _4303_ (.A1(_3153_),
    .A2(_0462_),
    .B1(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__a221oi_1 _4304_ (.A1(_0456_),
    .A2(_0455_),
    .B1(_0738_),
    .B2(_0459_),
    .C1(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__and4_1 _4305_ (.A(_0726_),
    .B(_0733_),
    .C(_0737_),
    .D(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__and2_1 _4306_ (.A(_0718_),
    .B(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__inv_2 _4307_ (.A(_0480_),
    .Y(_0744_));
 sky130_fd_sc_hd__clkbuf_4 _4308_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .X(_0745_));
 sky130_fd_sc_hd__nand2_1 _4309_ (.A(_0479_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__a22o_1 _4310_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_0747_));
 sky130_fd_sc_hd__inv_2 _4311_ (.A(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__o211a_1 _4312_ (.A1(_0744_),
    .A2(_0476_),
    .B1(_0746_),
    .C1(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__inv_2 _4313_ (.A(_0504_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_0503_),
    .B(_0520_),
    .Y(_0751_));
 sky130_fd_sc_hd__o21ai_1 _4315_ (.A1(_0750_),
    .A2(_0500_),
    .B1(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__a221oi_1 _4316_ (.A1(_0493_),
    .A2(_0492_),
    .B1(_0497_),
    .B2(_0496_),
    .C1(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_0514_),
    .B(_0508_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(_0519_),
    .B(_0522_),
    .Y(_0755_));
 sky130_fd_sc_hd__inv_2 _4319_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .Y(_0756_));
 sky130_fd_sc_hd__or2_1 _4320_ (.A(_0756_),
    .B(_0525_),
    .X(_0757_));
 sky130_fd_sc_hd__o2111a_1 _4321_ (.A1(_0472_),
    .A2(_0511_),
    .B1(_0754_),
    .C1(_0755_),
    .D1(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(_0538_),
    .B(_0528_),
    .Y(_0759_));
 sky130_fd_sc_hd__nand2_1 _4323_ (.A(_0543_),
    .B(_0539_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _4324_ (.A(_0759_),
    .B(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__a221oi_1 _4325_ (.A1(_0532_),
    .A2(_0531_),
    .B1(_0363_),
    .B2(_0535_),
    .C1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__and4_1 _4326_ (.A(_0749_),
    .B(_0753_),
    .C(_0758_),
    .D(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__inv_2 _4327_ (.A(_0558_),
    .Y(_0764_));
 sky130_fd_sc_hd__nand2_1 _4328_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_0765_));
 sky130_fd_sc_hd__nand2_1 _4329_ (.A(_0562_),
    .B(_0549_),
    .Y(_0766_));
 sky130_fd_sc_hd__inv_2 _4330_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0767_));
 sky130_fd_sc_hd__or2_1 _4331_ (.A(_0767_),
    .B(_0567_),
    .X(_0768_));
 sky130_fd_sc_hd__o2111a_1 _4332_ (.A1(_0764_),
    .A2(_0554_),
    .B1(_0765_),
    .C1(_0766_),
    .D1(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(_0575_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_0771_));
 sky130_fd_sc_hd__inv_2 _4335_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0772_));
 sky130_fd_sc_hd__or2_1 _4336_ (.A(_0772_),
    .B(_0583_),
    .X(_0773_));
 sky130_fd_sc_hd__o2111a_1 _4337_ (.A1(_0605_),
    .A2(_0572_),
    .B1(_0770_),
    .C1(_0771_),
    .D1(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__inv_2 _4338_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0775_));
 sky130_fd_sc_hd__or2_1 _4339_ (.A(_0775_),
    .B(_0596_),
    .X(_0776_));
 sky130_fd_sc_hd__o221a_1 _4340_ (.A1(_0594_),
    .A2(_0589_),
    .B1(_0587_),
    .B2(_0592_),
    .C1(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__inv_2 _4341_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_0778_));
 sky130_fd_sc_hd__o22ai_1 _4342_ (.A1(_0608_),
    .A2(_0607_),
    .B1(_0778_),
    .B2(_0610_),
    .Y(_0779_));
 sky130_fd_sc_hd__a221oi_1 _4343_ (.A1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .A2(_0601_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .B2(_0604_),
    .C1(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__and4_1 _4344_ (.A(_0769_),
    .B(_0774_),
    .C(_0777_),
    .D(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__and3_1 _4345_ (.A(_0743_),
    .B(_0763_),
    .C(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__buf_2 _4346_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0783_));
 sky130_fd_sc_hd__nand2_1 _4347_ (.A(_0618_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__nand3_1 _4348_ (.A(_0698_),
    .B(_0782_),
    .C(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__o21a_1 _4349_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .A2(_3043_),
    .B1(_2980_),
    .X(_0786_));
 sky130_fd_sc_hd__o21a_1 _4350_ (.A1(_3103_),
    .A2(_0785_),
    .B1(_0786_),
    .X(_0296_));
 sky130_fd_sc_hd__inv_2 _4351_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_0787_));
 sky130_fd_sc_hd__o22ai_1 _4352_ (.A1(_0623_),
    .A2(_3130_),
    .B1(_0787_),
    .B2(_3138_),
    .Y(_0788_));
 sky130_fd_sc_hd__a221oi_1 _4353_ (.A1(_3209_),
    .A2(_3115_),
    .B1(_3203_),
    .B2(_3122_),
    .C1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _4354_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_0790_));
 sky130_fd_sc_hd__nand2_1 _4355_ (.A(_3160_),
    .B(_3148_),
    .Y(_0791_));
 sky130_fd_sc_hd__o21ai_1 _4356_ (.A1(_0790_),
    .A2(_3156_),
    .B1(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__a221oi_1 _4357_ (.A1(_3175_),
    .A2(_3147_),
    .B1(_0630_),
    .B2(_3152_),
    .C1(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__nand2_1 _4358_ (.A(_3174_),
    .B(_3181_),
    .Y(_0794_));
 sky130_fd_sc_hd__buf_2 _4359_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(_3180_),
    .B(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__or2_1 _4361_ (.A(_3165_),
    .B(_3187_),
    .X(_0797_));
 sky130_fd_sc_hd__o2111a_1 _4362_ (.A1(_3132_),
    .A2(_3169_),
    .B1(_0794_),
    .C1(_0796_),
    .D1(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__clkbuf_4 _4363_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .X(_0799_));
 sky130_fd_sc_hd__nand2_1 _4364_ (.A(_3202_),
    .B(_3195_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(_3208_),
    .B(_3190_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(_0800_),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__a221oi_2 _4367_ (.A1(_0637_),
    .A2(_3194_),
    .B1(_0799_),
    .B2(_3198_),
    .C1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__and4_1 _4368_ (.A(_0789_),
    .B(_0793_),
    .C(_0798_),
    .D(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__inv_2 _4369_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_0805_));
 sky130_fd_sc_hd__o22ai_1 _4370_ (.A1(_0643_),
    .A2(_3224_),
    .B1(_0805_),
    .B2(_3227_),
    .Y(_0806_));
 sky130_fd_sc_hd__a221oi_1 _4371_ (.A1(_3078_),
    .A2(_3218_),
    .B1(_3081_),
    .B2(_3221_),
    .C1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__nand2_1 _4372_ (.A(_3241_),
    .B(_3090_),
    .Y(_0808_));
 sky130_fd_sc_hd__o21ai_1 _4373_ (.A1(_3269_),
    .A2(_3238_),
    .B1(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__a221oi_1 _4374_ (.A1(_3084_),
    .A2(_3232_),
    .B1(_3087_),
    .B2(_3235_),
    .C1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_2 _4375_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _4376_ (.A(_3256_),
    .B(_3062_),
    .Y(_0812_));
 sky130_fd_sc_hd__o21ai_1 _4377_ (.A1(_0811_),
    .A2(_3253_),
    .B1(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a221oi_1 _4378_ (.A1(_3065_),
    .A2(_3247_),
    .B1(_3068_),
    .B2(_3250_),
    .C1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _4379_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_0815_));
 sky130_fd_sc_hd__o22ai_1 _4380_ (.A1(_0653_),
    .A2(_3268_),
    .B1(_0815_),
    .B2(_3271_),
    .Y(_0816_));
 sky130_fd_sc_hd__a221oi_1 _4381_ (.A1(_0619_),
    .A2(_3262_),
    .B1(_0783_),
    .B2(_3265_),
    .C1(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__and4_1 _4382_ (.A(_0807_),
    .B(_0810_),
    .C(_0814_),
    .D(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__buf_2 _4383_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0819_));
 sky130_fd_sc_hd__inv_2 _4384_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_0820_));
 sky130_fd_sc_hd__o22ai_1 _4385_ (.A1(_0658_),
    .A2(_3288_),
    .B1(_0820_),
    .B2(_3291_),
    .Y(_0821_));
 sky130_fd_sc_hd__a221oi_1 _4386_ (.A1(_0657_),
    .A2(_3281_),
    .B1(_0819_),
    .B2(_3285_),
    .C1(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__nand2_1 _4387_ (.A(_3296_),
    .B(_3301_),
    .Y(_0823_));
 sky130_fd_sc_hd__clkbuf_4 _4388_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_0824_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_3300_),
    .B(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__nand2_1 _4390_ (.A(_3305_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0826_));
 sky130_fd_sc_hd__nand2_1 _4391_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0827_));
 sky130_fd_sc_hd__and4_1 _4392_ (.A(_0823_),
    .B(_0825_),
    .C(_0826_),
    .D(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__inv_2 _4393_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_0829_));
 sky130_fd_sc_hd__o22ai_1 _4394_ (.A1(_0668_),
    .A2(_3314_),
    .B1(_0829_),
    .B2(_3317_),
    .Y(_0830_));
 sky130_fd_sc_hd__clkbuf_4 _4395_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0831_));
 sky130_fd_sc_hd__a22o_1 _4396_ (.A1(_3320_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .B1(_3322_),
    .B2(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__nor2_1 _4397_ (.A(_0830_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_2 _4398_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_0834_));
 sky130_fd_sc_hd__o22ai_1 _4399_ (.A1(_0673_),
    .A2(_3336_),
    .B1(_0834_),
    .B2(_3339_),
    .Y(_0835_));
 sky130_fd_sc_hd__a221oi_1 _4400_ (.A1(_3366_),
    .A2(_3329_),
    .B1(_3370_),
    .B2(_3333_),
    .C1(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__and4_1 _4401_ (.A(_0822_),
    .B(_0828_),
    .C(_0833_),
    .D(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__nand2_1 _4402_ (.A(_3356_),
    .B(_3350_),
    .Y(_0838_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_3361_),
    .B(_3343_),
    .Y(_0839_));
 sky130_fd_sc_hd__nand2_1 _4404_ (.A(_0838_),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__a221oi_1 _4405_ (.A1(_3403_),
    .A2(_3349_),
    .B1(_3407_),
    .B2(_3353_),
    .C1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_3375_),
    .B(_0686_),
    .Y(_0842_));
 sky130_fd_sc_hd__nand2_1 _4407_ (.A(_3380_),
    .B(_3391_),
    .Y(_0843_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(_0842_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__a221oi_1 _4409_ (.A1(_3381_),
    .A2(_3369_),
    .B1(_3376_),
    .B2(_3372_),
    .C1(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__inv_2 _4410_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _4412_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0848_));
 sky130_fd_sc_hd__or2_1 _4413_ (.A(_3385_),
    .B(_3400_),
    .X(_0849_));
 sky130_fd_sc_hd__o2111a_1 _4414_ (.A1(_0846_),
    .A2(_3387_),
    .B1(_0847_),
    .C1(_0848_),
    .D1(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__buf_2 _4415_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_0852_));
 sky130_fd_sc_hd__o21ai_1 _4417_ (.A1(_0649_),
    .A2(_3413_),
    .B1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__a221oi_1 _4418_ (.A1(_0693_),
    .A2(_3406_),
    .B1(_0851_),
    .B2(_3410_),
    .C1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__and4_1 _4419_ (.A(_0841_),
    .B(_0845_),
    .C(_0850_),
    .D(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__and4_1 _4420_ (.A(_0804_),
    .B(_0818_),
    .C(_0837_),
    .D(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__nand2_1 _4421_ (.A(_0338_),
    .B(_0332_),
    .Y(_0857_));
 sky130_fd_sc_hd__nand2_1 _4422_ (.A(_0343_),
    .B(_0326_),
    .Y(_0858_));
 sky130_fd_sc_hd__nand2_1 _4423_ (.A(_0857_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__a221oi_1 _4424_ (.A1(_0381_),
    .A2(_0331_),
    .B1(_0385_),
    .B2(_0335_),
    .C1(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__inv_2 _4425_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_0861_));
 sky130_fd_sc_hd__o22ai_1 _4426_ (.A1(_0703_),
    .A2(_0350_),
    .B1(_0861_),
    .B2(_0353_),
    .Y(_0862_));
 sky130_fd_sc_hd__a22o_1 _4427_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .B1(_0359_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0863_));
 sky130_fd_sc_hd__nor2_1 _4428_ (.A(_0862_),
    .B(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__buf_2 _4429_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_0865_));
 sky130_fd_sc_hd__nand2_1 _4430_ (.A(_0376_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__o21ai_1 _4431_ (.A1(_0348_),
    .A2(_0373_),
    .B1(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__a221oi_1 _4432_ (.A1(_0707_),
    .A2(_0366_),
    .B1(_0377_),
    .B2(_0370_),
    .C1(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__buf_2 _4433_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_1 _4434_ (.A(_0394_),
    .B(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__o21ai_1 _4435_ (.A1(_0734_),
    .A2(_0391_),
    .B1(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__a221oi_1 _4436_ (.A1(_0713_),
    .A2(_0384_),
    .B1(_0714_),
    .B2(_0388_),
    .C1(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__and4_1 _4437_ (.A(_0860_),
    .B(_0864_),
    .C(_0868_),
    .D(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__buf_2 _4438_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _4439_ (.A(_0405_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__buf_2 _4440_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .X(_0876_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(_0409_),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__or2_1 _4442_ (.A(_0429_),
    .B(_0414_),
    .X(_0878_));
 sky130_fd_sc_hd__o2111a_1 _4443_ (.A1(_0412_),
    .A2(_0402_),
    .B1(_0875_),
    .C1(_0877_),
    .D1(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__inv_2 _4444_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _4445_ (.A(_0422_),
    .B(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0881_));
 sky130_fd_sc_hd__nand2_1 _4446_ (.A(_0426_),
    .B(_0452_),
    .Y(_0882_));
 sky130_fd_sc_hd__or2_1 _4447_ (.A(_0417_),
    .B(_0431_),
    .X(_0883_));
 sky130_fd_sc_hd__o2111a_1 _4448_ (.A1(_0880_),
    .A2(_0419_),
    .B1(_0881_),
    .C1(_0882_),
    .D1(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__inv_2 _4449_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_0885_));
 sky130_fd_sc_hd__nand2_1 _4450_ (.A(_0447_),
    .B(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_0886_));
 sky130_fd_sc_hd__o21ai_1 _4451_ (.A1(_0885_),
    .A2(_0444_),
    .B1(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__a221oi_1 _4452_ (.A1(_0410_),
    .A2(_0437_),
    .B1(_0722_),
    .B2(_0441_),
    .C1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__buf_2 _4453_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .X(_0889_));
 sky130_fd_sc_hd__buf_2 _4454_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .X(_0890_));
 sky130_fd_sc_hd__nand2_1 _4455_ (.A(_0465_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__o21ai_1 _4456_ (.A1(_0626_),
    .A2(_0462_),
    .B1(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__a221oi_1 _4457_ (.A1(_0738_),
    .A2(_0455_),
    .B1(_0889_),
    .B2(_0459_),
    .C1(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__and4_1 _4458_ (.A(_0879_),
    .B(_0884_),
    .C(_0888_),
    .D(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__and2_1 _4459_ (.A(_0873_),
    .B(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__inv_2 _4460_ (.A(_0745_),
    .Y(_0896_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_0479_),
    .B(_0486_),
    .Y(_0897_));
 sky130_fd_sc_hd__a22o_1 _4462_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_0898_));
 sky130_fd_sc_hd__inv_2 _4463_ (.A(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__o211a_1 _4464_ (.A1(_0896_),
    .A2(_0476_),
    .B1(_0897_),
    .C1(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__inv_2 _4465_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .Y(_0901_));
 sky130_fd_sc_hd__nand2_1 _4466_ (.A(_0503_),
    .B(_0522_),
    .Y(_0902_));
 sky130_fd_sc_hd__o21ai_1 _4467_ (.A1(_0901_),
    .A2(_0500_),
    .B1(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__a221oi_1 _4468_ (.A1(_0497_),
    .A2(_0492_),
    .B1(_0504_),
    .B2(_0496_),
    .C1(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__nand2_1 _4469_ (.A(_0514_),
    .B(_0471_),
    .Y(_0905_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_0519_),
    .B(_0515_),
    .Y(_0906_));
 sky130_fd_sc_hd__or2_1 _4471_ (.A(_0509_),
    .B(_0525_),
    .X(_0907_));
 sky130_fd_sc_hd__o2111a_1 _4472_ (.A1(_0744_),
    .A2(_0511_),
    .B1(_0905_),
    .C1(_0906_),
    .D1(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__nand2_1 _4473_ (.A(_0538_),
    .B(_0532_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_1 _4474_ (.A(_0543_),
    .B(_0528_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2_1 _4475_ (.A(_0909_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__a221oi_1 _4476_ (.A1(_0363_),
    .A2(_0531_),
    .B1(_0367_),
    .B2(_0535_),
    .C1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__and4_1 _4477_ (.A(_0900_),
    .B(_0904_),
    .C(_0908_),
    .D(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__nand2_1 _4478_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0914_));
 sky130_fd_sc_hd__nand2_1 _4479_ (.A(_0562_),
    .B(_0558_),
    .Y(_0915_));
 sky130_fd_sc_hd__or2_1 _4480_ (.A(_0581_),
    .B(_0567_),
    .X(_0916_));
 sky130_fd_sc_hd__o2111a_1 _4481_ (.A1(_0565_),
    .A2(_0554_),
    .B1(_0914_),
    .C1(_0915_),
    .D1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_0575_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0919_));
 sky130_fd_sc_hd__or2_1 _4484_ (.A(_0570_),
    .B(_0583_),
    .X(_0920_));
 sky130_fd_sc_hd__o2111a_1 _4485_ (.A1(_0608_),
    .A2(_0572_),
    .B1(_0918_),
    .C1(_0919_),
    .D1(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__or2_1 _4486_ (.A(_0550_),
    .B(_0596_),
    .X(_0922_));
 sky130_fd_sc_hd__o221a_1 _4487_ (.A1(_0775_),
    .A2(_0589_),
    .B1(_0594_),
    .B2(_0592_),
    .C1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__inv_2 _4488_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_0924_));
 sky130_fd_sc_hd__o22ai_1 _4489_ (.A1(_0778_),
    .A2(_0607_),
    .B1(_0924_),
    .B2(_0610_),
    .Y(_0925_));
 sky130_fd_sc_hd__a221oi_1 _4490_ (.A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .A2(_0601_),
    .B1(_0493_),
    .B2(_0604_),
    .C1(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__and4_1 _4491_ (.A(_0917_),
    .B(_0921_),
    .C(_0923_),
    .D(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__and3_1 _4492_ (.A(_0895_),
    .B(_0913_),
    .C(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(_0618_),
    .B(_0586_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand3_1 _4494_ (.A(_0856_),
    .B(_0928_),
    .C(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__inv_2 _4495_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_0931_));
 sky130_fd_sc_hd__buf_2 _4496_ (.A(_3102_),
    .X(_0932_));
 sky130_fd_sc_hd__a21oi_1 _4497_ (.A1(_0931_),
    .A2(_0932_),
    .B1(_2985_),
    .Y(_0933_));
 sky130_fd_sc_hd__o21a_1 _4498_ (.A1(_3103_),
    .A2(_0930_),
    .B1(_0933_),
    .X(_0295_));
 sky130_fd_sc_hd__inv_2 _4499_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_0934_));
 sky130_fd_sc_hd__o22ai_1 _4500_ (.A1(_0787_),
    .A2(_3130_),
    .B1(_0934_),
    .B2(_3138_),
    .Y(_0935_));
 sky130_fd_sc_hd__a221oi_1 _4501_ (.A1(_3203_),
    .A2(_3115_),
    .B1(_3190_),
    .B2(_3122_),
    .C1(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__inv_2 _4502_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _4503_ (.A(_3160_),
    .B(_3175_),
    .Y(_0938_));
 sky130_fd_sc_hd__o21ai_1 _4504_ (.A1(_0937_),
    .A2(_3156_),
    .B1(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__a221oi_1 _4505_ (.A1(_0630_),
    .A2(_3147_),
    .B1(_3181_),
    .B2(_3152_),
    .C1(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand2_1 _4506_ (.A(_3174_),
    .B(_0632_),
    .Y(_0941_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(_3180_),
    .B(_3131_),
    .Y(_0942_));
 sky130_fd_sc_hd__or2_1 _4508_ (.A(_3123_),
    .B(_3187_),
    .X(_0943_));
 sky130_fd_sc_hd__o2111a_1 _4509_ (.A1(_0623_),
    .A2(_3169_),
    .B1(_0941_),
    .C1(_0942_),
    .D1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__nand2_1 _4510_ (.A(_3202_),
    .B(_0637_),
    .Y(_0945_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_3208_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_0945_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__a221oi_2 _4513_ (.A1(_0799_),
    .A2(_3194_),
    .B1(_0661_),
    .B2(_3198_),
    .C1(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__and4_1 _4514_ (.A(_0936_),
    .B(_0940_),
    .C(_0944_),
    .D(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__inv_2 _4515_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_0950_));
 sky130_fd_sc_hd__o22ai_1 _4516_ (.A1(_0805_),
    .A2(_3224_),
    .B1(_0950_),
    .B2(_3227_),
    .Y(_0951_));
 sky130_fd_sc_hd__a221oi_1 _4517_ (.A1(_3081_),
    .A2(_3218_),
    .B1(_3084_),
    .B2(_3221_),
    .C1(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__nand2_1 _4518_ (.A(_3241_),
    .B(_3093_),
    .Y(_0953_));
 sky130_fd_sc_hd__o21ai_1 _4519_ (.A1(_0653_),
    .A2(_3238_),
    .B1(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__a221oi_1 _4520_ (.A1(_3087_),
    .A2(_3232_),
    .B1(_3090_),
    .B2(_3235_),
    .C1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__inv_2 _4521_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_0956_));
 sky130_fd_sc_hd__nand2_1 _4522_ (.A(_3256_),
    .B(_3065_),
    .Y(_0957_));
 sky130_fd_sc_hd__o21ai_1 _4523_ (.A1(_0956_),
    .A2(_3253_),
    .B1(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__a221oi_1 _4524_ (.A1(_3068_),
    .A2(_3247_),
    .B1(_3071_),
    .B2(_3250_),
    .C1(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_2 _4525_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_0960_));
 sky130_fd_sc_hd__o22ai_1 _4526_ (.A1(_0815_),
    .A2(_3268_),
    .B1(_0960_),
    .B2(_3271_),
    .Y(_0961_));
 sky130_fd_sc_hd__a221oi_1 _4527_ (.A1(_0783_),
    .A2(_3262_),
    .B1(_0586_),
    .B2(_3265_),
    .C1(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__and4_1 _4528_ (.A(_0952_),
    .B(_0955_),
    .C(_0959_),
    .D(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__o22ai_1 _4529_ (.A1(_0820_),
    .A2(_3288_),
    .B1(_3334_),
    .B2(_3291_),
    .Y(_0964_));
 sky130_fd_sc_hd__a221oi_1 _4530_ (.A1(_0819_),
    .A2(_3281_),
    .B1(_3326_),
    .B2(_3285_),
    .C1(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _4531_ (.A(_3296_),
    .B(_0663_),
    .Y(_0966_));
 sky130_fd_sc_hd__clkbuf_4 _4532_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_0967_));
 sky130_fd_sc_hd__nand2_1 _4533_ (.A(_3300_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_3305_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0969_));
 sky130_fd_sc_hd__nand2_1 _4535_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0970_));
 sky130_fd_sc_hd__and4_1 _4536_ (.A(_0966_),
    .B(_0968_),
    .C(_0969_),
    .D(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__o22ai_1 _4537_ (.A1(_0829_),
    .A2(_3314_),
    .B1(_3286_),
    .B2(_3317_),
    .Y(_0972_));
 sky130_fd_sc_hd__a22o_1 _4538_ (.A1(_3320_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .B1(_3322_),
    .B2(_3275_),
    .X(_0973_));
 sky130_fd_sc_hd__nor2_1 _4539_ (.A(_0972_),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__inv_2 _4540_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_0975_));
 sky130_fd_sc_hd__o22ai_1 _4541_ (.A1(_0834_),
    .A2(_3336_),
    .B1(_0975_),
    .B2(_3339_),
    .Y(_0976_));
 sky130_fd_sc_hd__a221oi_1 _4542_ (.A1(_3370_),
    .A2(_3329_),
    .B1(_3381_),
    .B2(_3333_),
    .C1(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__and4_1 _4543_ (.A(_0965_),
    .B(_0971_),
    .C(_0974_),
    .D(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__nand2_1 _4544_ (.A(_3356_),
    .B(_3403_),
    .Y(_0979_));
 sky130_fd_sc_hd__nand2_1 _4545_ (.A(_3361_),
    .B(_3350_),
    .Y(_0980_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(_0979_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__a221oi_1 _4547_ (.A1(_3407_),
    .A2(_3349_),
    .B1(_0693_),
    .B2(_3353_),
    .C1(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand2_1 _4548_ (.A(_3375_),
    .B(_3396_),
    .Y(_0983_));
 sky130_fd_sc_hd__nand2_1 _4549_ (.A(_3380_),
    .B(_0686_),
    .Y(_0984_));
 sky130_fd_sc_hd__nand2_1 _4550_ (.A(_0983_),
    .B(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__a221oi_1 _4551_ (.A1(_3376_),
    .A2(_3369_),
    .B1(_3391_),
    .B2(_3372_),
    .C1(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__inv_2 _4552_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_0987_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_0988_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_0989_));
 sky130_fd_sc_hd__or2_1 _4555_ (.A(_0685_),
    .B(_3400_),
    .X(_0990_));
 sky130_fd_sc_hd__o2111a_1 _4556_ (.A1(_0987_),
    .A2(_3387_),
    .B1(_0988_),
    .C1(_0989_),
    .D1(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_0992_));
 sky130_fd_sc_hd__o21ai_1 _4558_ (.A1(_0811_),
    .A2(_3413_),
    .B1(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__a221oi_1 _4559_ (.A1(_0851_),
    .A2(_3406_),
    .B1(_3044_),
    .B2(_3410_),
    .C1(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__and4_1 _4560_ (.A(_0982_),
    .B(_0986_),
    .C(_0991_),
    .D(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__and4_1 _4561_ (.A(_0949_),
    .B(_0963_),
    .C(_0978_),
    .D(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__nand2_1 _4562_ (.A(_0338_),
    .B(_0381_),
    .Y(_0997_));
 sky130_fd_sc_hd__nand2_1 _4563_ (.A(_0343_),
    .B(_0332_),
    .Y(_0998_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_0997_),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__a221oi_1 _4565_ (.A1(_0385_),
    .A2(_0331_),
    .B1(_0713_),
    .B2(_0335_),
    .C1(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__inv_2 _4566_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_1001_));
 sky130_fd_sc_hd__o22ai_1 _4567_ (.A1(_0861_),
    .A2(_0350_),
    .B1(_1001_),
    .B2(_0353_),
    .Y(_1002_));
 sky130_fd_sc_hd__a22o_1 _4568_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .B1(_0359_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_1003_));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(_1002_),
    .B(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand2_1 _4570_ (.A(_0376_),
    .B(_0357_),
    .Y(_1005_));
 sky130_fd_sc_hd__o21ai_1 _4571_ (.A1(_0351_),
    .A2(_0373_),
    .B1(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__a221oi_1 _4572_ (.A1(_0377_),
    .A2(_0366_),
    .B1(_0709_),
    .B2(_0370_),
    .C1(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__nand2_1 _4573_ (.A(_0394_),
    .B(_0448_),
    .Y(_1008_));
 sky130_fd_sc_hd__o21ai_1 _4574_ (.A1(_0885_),
    .A2(_0391_),
    .B1(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__a221oi_1 _4575_ (.A1(_0714_),
    .A2(_0384_),
    .B1(_0869_),
    .B2(_0388_),
    .C1(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__and4_1 _4576_ (.A(_1000_),
    .B(_1004_),
    .C(_1007_),
    .D(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_4 _4577_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .X(_1012_));
 sky130_fd_sc_hd__nand2_1 _4578_ (.A(_0405_),
    .B(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__nand2_1 _4579_ (.A(_0409_),
    .B(_0720_),
    .Y(_1014_));
 sky130_fd_sc_hd__or2_1 _4580_ (.A(_0731_),
    .B(_0414_),
    .X(_1015_));
 sky130_fd_sc_hd__o2111a_1 _4581_ (.A1(_0724_),
    .A2(_0402_),
    .B1(_1013_),
    .C1(_1014_),
    .D1(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__inv_2 _4582_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_1017_));
 sky130_fd_sc_hd__nand2_1 _4583_ (.A(_0422_),
    .B(_0729_),
    .Y(_1018_));
 sky130_fd_sc_hd__nand2_1 _4584_ (.A(_0426_),
    .B(_0456_),
    .Y(_1019_));
 sky130_fd_sc_hd__or2_1 _4585_ (.A(_0727_),
    .B(_0431_),
    .X(_1020_));
 sky130_fd_sc_hd__o2111a_1 _4586_ (.A1(_1017_),
    .A2(_0419_),
    .B1(_1018_),
    .C1(_1019_),
    .D1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__inv_2 _4587_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2_1 _4588_ (.A(_0447_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1023_));
 sky130_fd_sc_hd__o21ai_1 _4589_ (.A1(_1022_),
    .A2(_0444_),
    .B1(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__a221oi_1 _4590_ (.A1(_0722_),
    .A2(_0437_),
    .B1(_0876_),
    .B2(_0441_),
    .C1(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(_0465_),
    .B(_3161_),
    .Y(_1026_));
 sky130_fd_sc_hd__o21ai_1 _4592_ (.A1(_0790_),
    .A2(_0462_),
    .B1(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__a221oi_1 _4593_ (.A1(_0889_),
    .A2(_0455_),
    .B1(_0890_),
    .B2(_0459_),
    .C1(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__and4_1 _4594_ (.A(_1016_),
    .B(_1021_),
    .C(_1025_),
    .D(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__and2_1 _4595_ (.A(_1011_),
    .B(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__inv_2 _4596_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_1031_));
 sky130_fd_sc_hd__nand2_1 _4597_ (.A(_0479_),
    .B(_0544_),
    .Y(_1032_));
 sky130_fd_sc_hd__a22o_1 _4598_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_1033_));
 sky130_fd_sc_hd__inv_2 _4599_ (.A(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__o211a_1 _4600_ (.A1(_1031_),
    .A2(_0476_),
    .B1(_1032_),
    .C1(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__nand2_1 _4601_ (.A(_0503_),
    .B(_0515_),
    .Y(_1036_));
 sky130_fd_sc_hd__o21ai_1 _4602_ (.A1(_0523_),
    .A2(_0500_),
    .B1(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__a221oi_1 _4603_ (.A1(_0504_),
    .A2(_0492_),
    .B1(_0520_),
    .B2(_0496_),
    .C1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__nand2_1 _4604_ (.A(_0514_),
    .B(_0480_),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _4605_ (.A(_0519_),
    .B(_0508_),
    .Y(_1040_));
 sky130_fd_sc_hd__or2_1 _4606_ (.A(_0472_),
    .B(_0525_),
    .X(_1041_));
 sky130_fd_sc_hd__o2111a_1 _4607_ (.A1(_0896_),
    .A2(_0511_),
    .B1(_1039_),
    .C1(_1040_),
    .D1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__nand2_1 _4608_ (.A(_0538_),
    .B(_0363_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _4609_ (.A(_0543_),
    .B(_0532_),
    .Y(_1044_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(_1043_),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a221oi_1 _4611_ (.A1(_0367_),
    .A2(_0531_),
    .B1(_0707_),
    .B2(_0535_),
    .C1(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__and4_1 _4612_ (.A(_1035_),
    .B(_1038_),
    .C(_1042_),
    .D(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__nand2_1 _4613_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_1 _4614_ (.A(_0562_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_1049_));
 sky130_fd_sc_hd__or2_1 _4615_ (.A(_0772_),
    .B(_0567_),
    .X(_1050_));
 sky130_fd_sc_hd__o2111a_1 _4616_ (.A1(_0767_),
    .A2(_0554_),
    .B1(_1048_),
    .C1(_1049_),
    .D1(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__nand2_1 _4617_ (.A(_0575_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _4618_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1053_));
 sky130_fd_sc_hd__or2_1 _4619_ (.A(_0605_),
    .B(_0583_),
    .X(_1054_));
 sky130_fd_sc_hd__o2111a_1 _4620_ (.A1(_0778_),
    .A2(_0572_),
    .B1(_1052_),
    .C1(_1053_),
    .D1(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__or2_1 _4621_ (.A(_0764_),
    .B(_0596_),
    .X(_1056_));
 sky130_fd_sc_hd__o221a_1 _4622_ (.A1(_0550_),
    .A2(_0589_),
    .B1(_0775_),
    .B2(_0592_),
    .C1(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__inv_2 _4623_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1058_));
 sky130_fd_sc_hd__o22ai_1 _4624_ (.A1(_0924_),
    .A2(_0607_),
    .B1(_1058_),
    .B2(_0610_),
    .Y(_1059_));
 sky130_fd_sc_hd__a221oi_1 _4625_ (.A1(_0493_),
    .A2(_0601_),
    .B1(_0497_),
    .B2(_0604_),
    .C1(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__and4_1 _4626_ (.A(_1051_),
    .B(_1055_),
    .C(_1057_),
    .D(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__and3_1 _4627_ (.A(_1030_),
    .B(_1047_),
    .C(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__nand2_1 _4628_ (.A(_0618_),
    .B(_0593_),
    .Y(_1063_));
 sky130_fd_sc_hd__nand3_1 _4629_ (.A(_0996_),
    .B(_1062_),
    .C(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__inv_2 _4630_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_1065_));
 sky130_fd_sc_hd__a21oi_1 _4631_ (.A1(_1065_),
    .A2(_0932_),
    .B1(_2985_),
    .Y(_1066_));
 sky130_fd_sc_hd__o21a_1 _4632_ (.A1(_3103_),
    .A2(_1064_),
    .B1(_1066_),
    .X(_0294_));
 sky130_fd_sc_hd__inv_2 _4633_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1067_));
 sky130_fd_sc_hd__o22ai_1 _4634_ (.A1(_0934_),
    .A2(_3130_),
    .B1(_1067_),
    .B2(_3138_),
    .Y(_1068_));
 sky130_fd_sc_hd__a221oi_1 _4635_ (.A1(_3190_),
    .A2(_3115_),
    .B1(_3195_),
    .B2(_3122_),
    .C1(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__inv_2 _4636_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1070_));
 sky130_fd_sc_hd__nand2_1 _4637_ (.A(_3160_),
    .B(_0630_),
    .Y(_1071_));
 sky130_fd_sc_hd__o21ai_1 _4638_ (.A1(_1070_),
    .A2(_3156_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__a221oi_1 _4639_ (.A1(_3181_),
    .A2(_3147_),
    .B1(_0632_),
    .B2(_3152_),
    .C1(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__nand2_1 _4640_ (.A(_3174_),
    .B(_0795_),
    .Y(_1074_));
 sky130_fd_sc_hd__nand2_1 _4641_ (.A(_3180_),
    .B(_3104_),
    .Y(_1075_));
 sky130_fd_sc_hd__or2_1 _4642_ (.A(_3132_),
    .B(_3187_),
    .X(_1076_));
 sky130_fd_sc_hd__o2111a_1 _4643_ (.A1(_0787_),
    .A2(_3169_),
    .B1(_1074_),
    .C1(_1075_),
    .D1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_1 _4644_ (.A(_3202_),
    .B(_0799_),
    .Y(_1078_));
 sky130_fd_sc_hd__nand2_1 _4645_ (.A(_3208_),
    .B(_0637_),
    .Y(_1079_));
 sky130_fd_sc_hd__nand2_1 _4646_ (.A(_1078_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__a221oi_2 _4647_ (.A1(_0661_),
    .A2(_3194_),
    .B1(_3301_),
    .B2(_3198_),
    .C1(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__and4_1 _4648_ (.A(_1069_),
    .B(_1073_),
    .C(_1077_),
    .D(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__inv_2 _4649_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1083_));
 sky130_fd_sc_hd__o22ai_1 _4650_ (.A1(_0950_),
    .A2(_3224_),
    .B1(_1083_),
    .B2(_3227_),
    .Y(_1084_));
 sky130_fd_sc_hd__a221oi_1 _4651_ (.A1(_3084_),
    .A2(_3218_),
    .B1(_3087_),
    .B2(_3221_),
    .C1(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__nand2_1 _4652_ (.A(_3241_),
    .B(_3096_),
    .Y(_1086_));
 sky130_fd_sc_hd__o21ai_1 _4653_ (.A1(_0815_),
    .A2(_3238_),
    .B1(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__a221oi_1 _4654_ (.A1(_3090_),
    .A2(_3232_),
    .B1(_3093_),
    .B2(_3235_),
    .C1(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__nand2_1 _4655_ (.A(_3256_),
    .B(_3068_),
    .Y(_1089_));
 sky130_fd_sc_hd__o21ai_1 _4656_ (.A1(_3222_),
    .A2(_3253_),
    .B1(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__a221oi_1 _4657_ (.A1(_3071_),
    .A2(_3247_),
    .B1(_3074_),
    .B2(_3250_),
    .C1(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__o22ai_1 _4658_ (.A1(_0960_),
    .A2(_3268_),
    .B1(_0590_),
    .B2(_3271_),
    .Y(_1092_));
 sky130_fd_sc_hd__a221oi_1 _4659_ (.A1(_0586_),
    .A2(_3262_),
    .B1(_0593_),
    .B2(_3265_),
    .C1(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__and4_1 _4660_ (.A(_1085_),
    .B(_1088_),
    .C(_1091_),
    .D(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__o22ai_1 _4661_ (.A1(_3334_),
    .A2(_3288_),
    .B1(_3337_),
    .B2(_3291_),
    .Y(_1095_));
 sky130_fd_sc_hd__a221oi_1 _4662_ (.A1(_3326_),
    .A2(_3281_),
    .B1(_3330_),
    .B2(_3285_),
    .C1(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_3296_),
    .B(_0824_),
    .Y(_1097_));
 sky130_fd_sc_hd__nand2_1 _4664_ (.A(_3300_),
    .B(_3323_),
    .Y(_1098_));
 sky130_fd_sc_hd__nand2_1 _4665_ (.A(_3305_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_1099_));
 sky130_fd_sc_hd__nand2_1 _4666_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_1100_));
 sky130_fd_sc_hd__and4_1 _4667_ (.A(_1097_),
    .B(_1098_),
    .C(_1099_),
    .D(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__o22ai_1 _4668_ (.A1(_3286_),
    .A2(_3314_),
    .B1(_3289_),
    .B2(_3317_),
    .Y(_1102_));
 sky130_fd_sc_hd__a22o_1 _4669_ (.A1(_3320_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .B1(_3322_),
    .B2(_3282_),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_1 _4670_ (.A(_1102_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__inv_2 _4671_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_1105_));
 sky130_fd_sc_hd__o22ai_1 _4672_ (.A1(_0975_),
    .A2(_3336_),
    .B1(_1105_),
    .B2(_3339_),
    .Y(_1106_));
 sky130_fd_sc_hd__a221oi_1 _4673_ (.A1(_3381_),
    .A2(_3329_),
    .B1(_3376_),
    .B2(_3333_),
    .C1(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__and4_1 _4674_ (.A(_1096_),
    .B(_1101_),
    .C(_1104_),
    .D(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__nand2_1 _4675_ (.A(_3356_),
    .B(_3407_),
    .Y(_1109_));
 sky130_fd_sc_hd__nand2_1 _4676_ (.A(_3361_),
    .B(_3403_),
    .Y(_1110_));
 sky130_fd_sc_hd__nand2_1 _4677_ (.A(_1109_),
    .B(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__a221oi_1 _4678_ (.A1(_0693_),
    .A2(_3349_),
    .B1(_0851_),
    .B2(_3353_),
    .C1(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_1 _4679_ (.A(_3375_),
    .B(_0688_),
    .Y(_1113_));
 sky130_fd_sc_hd__nand2_1 _4680_ (.A(_3380_),
    .B(_3396_),
    .Y(_1114_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_1113_),
    .B(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__a221oi_1 _4682_ (.A1(_3391_),
    .A2(_3369_),
    .B1(_0686_),
    .B2(_3372_),
    .C1(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__inv_2 _4683_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2_1 _4684_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_1118_));
 sky130_fd_sc_hd__nand2_1 _4685_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1119_));
 sky130_fd_sc_hd__or2_1 _4686_ (.A(_0846_),
    .B(_3400_),
    .X(_1120_));
 sky130_fd_sc_hd__o2111a_1 _4687_ (.A1(_1117_),
    .A2(_3387_),
    .B1(_1118_),
    .C1(_1119_),
    .D1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_1122_));
 sky130_fd_sc_hd__o21ai_1 _4689_ (.A1(_0956_),
    .A2(_3413_),
    .B1(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__a221oi_1 _4690_ (.A1(_3044_),
    .A2(_3406_),
    .B1(_3056_),
    .B2(_3410_),
    .C1(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__and4_1 _4691_ (.A(_1112_),
    .B(_1116_),
    .C(_1121_),
    .D(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__and4_1 _4692_ (.A(_1082_),
    .B(_1094_),
    .C(_1108_),
    .D(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__nand2_1 _4693_ (.A(_0338_),
    .B(_0385_),
    .Y(_1127_));
 sky130_fd_sc_hd__nand2_1 _4694_ (.A(_0343_),
    .B(_0381_),
    .Y(_1128_));
 sky130_fd_sc_hd__nand2_1 _4695_ (.A(_1127_),
    .B(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__a221oi_1 _4696_ (.A1(_0713_),
    .A2(_0331_),
    .B1(_0714_),
    .B2(_0335_),
    .C1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__inv_2 _4697_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_1131_));
 sky130_fd_sc_hd__o22ai_1 _4698_ (.A1(_1001_),
    .A2(_0350_),
    .B1(_1131_),
    .B2(_0353_),
    .Y(_1132_));
 sky130_fd_sc_hd__a22o_1 _4699_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .B1(_0359_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_1133_));
 sky130_fd_sc_hd__nor2_1 _4700_ (.A(_1132_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__nand2_1 _4701_ (.A(_0376_),
    .B(_0360_),
    .Y(_1135_));
 sky130_fd_sc_hd__o21ai_1 _4702_ (.A1(_0703_),
    .A2(_0373_),
    .B1(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__a221oi_1 _4703_ (.A1(_0709_),
    .A2(_0366_),
    .B1(_0865_),
    .B2(_0370_),
    .C1(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__nand2_1 _4704_ (.A(_0394_),
    .B(_0434_),
    .Y(_1138_));
 sky130_fd_sc_hd__o21ai_1 _4705_ (.A1(_1022_),
    .A2(_0391_),
    .B1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__a221oi_1 _4706_ (.A1(_0869_),
    .A2(_0384_),
    .B1(_0448_),
    .B2(_0388_),
    .C1(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__and4_1 _4707_ (.A(_1130_),
    .B(_1134_),
    .C(_1137_),
    .D(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__nand2_1 _4708_ (.A(_0405_),
    .B(_0427_),
    .Y(_1142_));
 sky130_fd_sc_hd__nand2_1 _4709_ (.A(_0409_),
    .B(_0874_),
    .Y(_1143_));
 sky130_fd_sc_hd__or2_1 _4710_ (.A(_0417_),
    .B(_0414_),
    .X(_1144_));
 sky130_fd_sc_hd__o2111a_1 _4711_ (.A1(_0429_),
    .A2(_0402_),
    .B1(_1142_),
    .C1(_1143_),
    .D1(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__nand2_1 _4712_ (.A(_0422_),
    .B(_0452_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _4713_ (.A(_0426_),
    .B(_0738_),
    .Y(_1147_));
 sky130_fd_sc_hd__or2_1 _4714_ (.A(_0880_),
    .B(_0431_),
    .X(_1148_));
 sky130_fd_sc_hd__o2111a_1 _4715_ (.A1(_0460_),
    .A2(_0419_),
    .B1(_1146_),
    .C1(_1147_),
    .D1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__inv_2 _4716_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_1 _4717_ (.A(_0447_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1151_));
 sky130_fd_sc_hd__o21ai_1 _4718_ (.A1(_1150_),
    .A2(_0444_),
    .B1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__a221oi_1 _4719_ (.A1(_0876_),
    .A2(_0437_),
    .B1(_0720_),
    .B2(_0441_),
    .C1(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_1 _4720_ (.A(_0465_),
    .B(_3141_),
    .Y(_1154_));
 sky130_fd_sc_hd__o21ai_1 _4721_ (.A1(_0937_),
    .A2(_0462_),
    .B1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__a221oi_1 _4722_ (.A1(_0890_),
    .A2(_0455_),
    .B1(_3161_),
    .B2(_0459_),
    .C1(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__and4_1 _4723_ (.A(_1145_),
    .B(_1149_),
    .C(_1153_),
    .D(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__and2_1 _4724_ (.A(_1141_),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__inv_2 _4725_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_1 _4726_ (.A(_0479_),
    .B(_0539_),
    .Y(_1160_));
 sky130_fd_sc_hd__a22o_1 _4727_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_1161_));
 sky130_fd_sc_hd__inv_2 _4728_ (.A(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__o211a_1 _4729_ (.A1(_1159_),
    .A2(_0476_),
    .B1(_1160_),
    .C1(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(_0503_),
    .B(_0508_),
    .Y(_1164_));
 sky130_fd_sc_hd__o21ai_1 _4731_ (.A1(_0756_),
    .A2(_0500_),
    .B1(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a221oi_1 _4732_ (.A1(_0520_),
    .A2(_0492_),
    .B1(_0522_),
    .B2(_0496_),
    .C1(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_0514_),
    .B(_0745_),
    .Y(_1167_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(_0519_),
    .B(_0471_),
    .Y(_1168_));
 sky130_fd_sc_hd__or2_1 _4735_ (.A(_0744_),
    .B(_0525_),
    .X(_1169_));
 sky130_fd_sc_hd__o2111a_1 _4736_ (.A1(_1031_),
    .A2(_0511_),
    .B1(_1167_),
    .C1(_1168_),
    .D1(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nand2_1 _4737_ (.A(_0538_),
    .B(_0367_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0543_),
    .B(_0363_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(_1171_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__a221oi_1 _4740_ (.A1(_0707_),
    .A2(_0531_),
    .B1(_0377_),
    .B2(_0535_),
    .C1(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__and4_1 _4741_ (.A(_1163_),
    .B(_1166_),
    .C(_1170_),
    .D(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__nand2_1 _4742_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _4743_ (.A(_0562_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_1177_));
 sky130_fd_sc_hd__or2_1 _4744_ (.A(_0570_),
    .B(_0567_),
    .X(_1178_));
 sky130_fd_sc_hd__o2111a_1 _4745_ (.A1(_0581_),
    .A2(_0554_),
    .B1(_1176_),
    .C1(_1177_),
    .D1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__nand2_1 _4746_ (.A(_0575_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1180_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1181_));
 sky130_fd_sc_hd__or2_1 _4748_ (.A(_0608_),
    .B(_0583_),
    .X(_1182_));
 sky130_fd_sc_hd__o2111a_1 _4749_ (.A1(_0924_),
    .A2(_0572_),
    .B1(_1180_),
    .C1(_1181_),
    .D1(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__or2_1 _4750_ (.A(_0565_),
    .B(_0596_),
    .X(_1184_));
 sky130_fd_sc_hd__o221a_1 _4751_ (.A1(_0764_),
    .A2(_0589_),
    .B1(_0550_),
    .B2(_0592_),
    .C1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__inv_2 _4752_ (.A(_0493_),
    .Y(_1186_));
 sky130_fd_sc_hd__o22ai_1 _4753_ (.A1(_1058_),
    .A2(_0607_),
    .B1(_1186_),
    .B2(_0610_),
    .Y(_1187_));
 sky130_fd_sc_hd__a221oi_1 _4754_ (.A1(_0497_),
    .A2(_0601_),
    .B1(_0504_),
    .B2(_0604_),
    .C1(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__and4_1 _4755_ (.A(_1179_),
    .B(_1183_),
    .C(_1185_),
    .D(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__and3_1 _4756_ (.A(_1158_),
    .B(_1175_),
    .C(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_0618_),
    .B(_0563_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand3_1 _4758_ (.A(_1126_),
    .B(_1190_),
    .C(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__inv_4 _4759_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_1193_));
 sky130_fd_sc_hd__a21oi_1 _4760_ (.A1(_1193_),
    .A2(_0932_),
    .B1(_2985_),
    .Y(_1194_));
 sky130_fd_sc_hd__o21a_1 _4761_ (.A1(_3103_),
    .A2(_1192_),
    .B1(_1194_),
    .X(_0293_));
 sky130_fd_sc_hd__inv_2 _4762_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1195_));
 sky130_fd_sc_hd__o22ai_1 _4763_ (.A1(_1067_),
    .A2(_3130_),
    .B1(_1195_),
    .B2(_3138_),
    .Y(_1196_));
 sky130_fd_sc_hd__a221oi_1 _4764_ (.A1(_3195_),
    .A2(_3115_),
    .B1(_0637_),
    .B2(_3122_),
    .C1(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_1 _4765_ (.A(_3160_),
    .B(_3181_),
    .Y(_1198_));
 sky130_fd_sc_hd__o21ai_1 _4766_ (.A1(_3183_),
    .A2(_3156_),
    .B1(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__a221oi_1 _4767_ (.A1(_0632_),
    .A2(_3147_),
    .B1(_0795_),
    .B2(_3152_),
    .C1(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_3174_),
    .B(_3131_),
    .Y(_1201_));
 sky130_fd_sc_hd__nand2_1 _4769_ (.A(_3180_),
    .B(_3116_),
    .Y(_1202_));
 sky130_fd_sc_hd__or2_1 _4770_ (.A(_0623_),
    .B(_3187_),
    .X(_1203_));
 sky130_fd_sc_hd__o2111a_1 _4771_ (.A1(_0934_),
    .A2(_3169_),
    .B1(_1201_),
    .C1(_1202_),
    .D1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__nand2_1 _4772_ (.A(_3202_),
    .B(_0661_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand2_1 _4773_ (.A(_3208_),
    .B(_0799_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__a221oi_2 _4775_ (.A1(_3301_),
    .A2(_3194_),
    .B1(_0663_),
    .B2(_3198_),
    .C1(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__and4_1 _4776_ (.A(_1197_),
    .B(_1200_),
    .C(_1204_),
    .D(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__inv_2 _4777_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1210_));
 sky130_fd_sc_hd__o22ai_1 _4778_ (.A1(_1083_),
    .A2(_3224_),
    .B1(_1210_),
    .B2(_3227_),
    .Y(_1211_));
 sky130_fd_sc_hd__a221oi_1 _4779_ (.A1(_3087_),
    .A2(_3218_),
    .B1(_3090_),
    .B2(_3221_),
    .C1(_1211_),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _4780_ (.A(_3241_),
    .B(_3099_),
    .Y(_1213_));
 sky130_fd_sc_hd__o21ai_1 _4781_ (.A1(_0960_),
    .A2(_3238_),
    .B1(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__a221oi_1 _4782_ (.A1(_3093_),
    .A2(_3232_),
    .B1(_3096_),
    .B2(_3235_),
    .C1(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_1 _4783_ (.A(_3256_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1216_));
 sky130_fd_sc_hd__o21ai_1 _4784_ (.A1(_3225_),
    .A2(_3253_),
    .B1(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__a221oi_1 _4785_ (.A1(_3074_),
    .A2(_3247_),
    .B1(_3078_),
    .B2(_3250_),
    .C1(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__o22ai_1 _4786_ (.A1(_0590_),
    .A2(_3268_),
    .B1(_0587_),
    .B2(_3271_),
    .Y(_1219_));
 sky130_fd_sc_hd__a221oi_2 _4787_ (.A1(_0593_),
    .A2(_3262_),
    .B1(_0563_),
    .B2(_3265_),
    .C1(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__and4_1 _4788_ (.A(_1212_),
    .B(_1215_),
    .C(_1218_),
    .D(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__o22ai_1 _4789_ (.A1(_3337_),
    .A2(_3288_),
    .B1(_0673_),
    .B2(_3291_),
    .Y(_1222_));
 sky130_fd_sc_hd__a221oi_1 _4790_ (.A1(_3330_),
    .A2(_3281_),
    .B1(_3366_),
    .B2(_3285_),
    .C1(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_1 _4791_ (.A(_3296_),
    .B(_0967_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2_1 _4792_ (.A(_3300_),
    .B(_0670_),
    .Y(_1225_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_3305_),
    .B(_0824_),
    .Y(_1226_));
 sky130_fd_sc_hd__nand2_1 _4794_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1227_));
 sky130_fd_sc_hd__and4_1 _4795_ (.A(_1224_),
    .B(_1225_),
    .C(_1226_),
    .D(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__o22ai_1 _4796_ (.A1(_3289_),
    .A2(_3314_),
    .B1(_0658_),
    .B2(_3317_),
    .Y(_1229_));
 sky130_fd_sc_hd__a22o_1 _4797_ (.A1(_3320_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .B1(_3322_),
    .B2(_0657_),
    .X(_1230_));
 sky130_fd_sc_hd__nor2_1 _4798_ (.A(_1229_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__inv_2 _4799_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .Y(_1232_));
 sky130_fd_sc_hd__o22ai_1 _4800_ (.A1(_1105_),
    .A2(_3336_),
    .B1(_1232_),
    .B2(_3339_),
    .Y(_1233_));
 sky130_fd_sc_hd__a221oi_1 _4801_ (.A1(_3376_),
    .A2(_3329_),
    .B1(_3391_),
    .B2(_3333_),
    .C1(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__and4_1 _4802_ (.A(_1223_),
    .B(_1228_),
    .C(_1231_),
    .D(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__nand2_1 _4803_ (.A(_3356_),
    .B(_0693_),
    .Y(_1236_));
 sky130_fd_sc_hd__nand2_1 _4804_ (.A(_3361_),
    .B(_3407_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _4805_ (.A(_1236_),
    .B(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__a221oi_1 _4806_ (.A1(_0851_),
    .A2(_3349_),
    .B1(_3044_),
    .B2(_3353_),
    .C1(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(_3375_),
    .B(_3362_),
    .Y(_1240_));
 sky130_fd_sc_hd__nand2_1 _4808_ (.A(_3380_),
    .B(_0688_),
    .Y(_1241_));
 sky130_fd_sc_hd__nand2_1 _4809_ (.A(_1240_),
    .B(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__a221oi_1 _4810_ (.A1(_0686_),
    .A2(_3369_),
    .B1(_3396_),
    .B2(_3372_),
    .C1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__inv_2 _4811_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1244_));
 sky130_fd_sc_hd__nand2_1 _4812_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_1245_));
 sky130_fd_sc_hd__nand2_1 _4813_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1246_));
 sky130_fd_sc_hd__or2_1 _4814_ (.A(_0987_),
    .B(_3400_),
    .X(_1247_));
 sky130_fd_sc_hd__o2111a_1 _4815_ (.A1(_1244_),
    .A2(_3387_),
    .B1(_1245_),
    .C1(_1246_),
    .D1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__nand2_1 _4816_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_1249_));
 sky130_fd_sc_hd__o21ai_1 _4817_ (.A1(_3222_),
    .A2(_3413_),
    .B1(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__a221oi_1 _4818_ (.A1(_3056_),
    .A2(_3406_),
    .B1(_3059_),
    .B2(_3410_),
    .C1(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__and4_1 _4819_ (.A(_1239_),
    .B(_1243_),
    .C(_1248_),
    .D(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__and4_1 _4820_ (.A(_1209_),
    .B(_1221_),
    .C(_1235_),
    .D(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(_0338_),
    .B(_0713_),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _4822_ (.A(_0343_),
    .B(_0385_),
    .Y(_1255_));
 sky130_fd_sc_hd__nand2_1 _4823_ (.A(_1254_),
    .B(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__a221oi_1 _4824_ (.A1(_0714_),
    .A2(_0331_),
    .B1(_0869_),
    .B2(_0335_),
    .C1(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__inv_2 _4825_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1258_));
 sky130_fd_sc_hd__o22ai_1 _4826_ (.A1(_1131_),
    .A2(_0350_),
    .B1(_1258_),
    .B2(_0353_),
    .Y(_1259_));
 sky130_fd_sc_hd__a22o_1 _4827_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .B1(_0359_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_1260_));
 sky130_fd_sc_hd__nor2_1 _4828_ (.A(_1259_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand2_1 _4829_ (.A(_0376_),
    .B(_0344_),
    .Y(_1262_));
 sky130_fd_sc_hd__o21ai_1 _4830_ (.A1(_0861_),
    .A2(_0373_),
    .B1(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__a221oi_1 _4831_ (.A1(_0865_),
    .A2(_0366_),
    .B1(_0357_),
    .B2(_0370_),
    .C1(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_0394_),
    .B(_0438_),
    .Y(_1265_));
 sky130_fd_sc_hd__o21ai_1 _4833_ (.A1(_1150_),
    .A2(_0391_),
    .B1(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__a221oi_1 _4834_ (.A1(_0448_),
    .A2(_0384_),
    .B1(_0434_),
    .B2(_0388_),
    .C1(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__and4_1 _4835_ (.A(_1257_),
    .B(_1261_),
    .C(_1264_),
    .D(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__nand2_1 _4836_ (.A(_0405_),
    .B(_0729_),
    .Y(_1269_));
 sky130_fd_sc_hd__nand2_1 _4837_ (.A(_0409_),
    .B(_1012_),
    .Y(_1270_));
 sky130_fd_sc_hd__or2_1 _4838_ (.A(_0727_),
    .B(_0414_),
    .X(_1271_));
 sky130_fd_sc_hd__o2111a_1 _4839_ (.A1(_0731_),
    .A2(_0402_),
    .B1(_1269_),
    .C1(_1270_),
    .D1(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__nand2_1 _4840_ (.A(_0422_),
    .B(_0456_),
    .Y(_1273_));
 sky130_fd_sc_hd__nand2_1 _4841_ (.A(_0426_),
    .B(_0889_),
    .Y(_1274_));
 sky130_fd_sc_hd__or2_1 _4842_ (.A(_1017_),
    .B(_0431_),
    .X(_1275_));
 sky130_fd_sc_hd__o2111a_1 _4843_ (.A1(_3153_),
    .A2(_0419_),
    .B1(_1273_),
    .C1(_1274_),
    .D1(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(_0447_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1277_));
 sky130_fd_sc_hd__o21ai_1 _4845_ (.A1(_0399_),
    .A2(_0444_),
    .B1(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__a221oi_1 _4846_ (.A1(_0720_),
    .A2(_0437_),
    .B1(_0874_),
    .B2(_0441_),
    .C1(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(_0465_),
    .B(_3148_),
    .Y(_1280_));
 sky130_fd_sc_hd__o21ai_1 _4848_ (.A1(_1070_),
    .A2(_0462_),
    .B1(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__a221oi_1 _4849_ (.A1(_3161_),
    .A2(_0455_),
    .B1(_3141_),
    .B2(_0459_),
    .C1(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__and4_1 _4850_ (.A(_1272_),
    .B(_1276_),
    .C(_1279_),
    .D(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__and2_1 _4851_ (.A(_1268_),
    .B(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__inv_2 _4852_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_1285_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_0479_),
    .B(_0528_),
    .Y(_1286_));
 sky130_fd_sc_hd__a22o_1 _4854_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_1287_));
 sky130_fd_sc_hd__inv_2 _4855_ (.A(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hd__o211a_1 _4856_ (.A1(_1285_),
    .A2(_0476_),
    .B1(_1286_),
    .C1(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(_0503_),
    .B(_0471_),
    .Y(_1290_));
 sky130_fd_sc_hd__o21ai_1 _4858_ (.A1(_0509_),
    .A2(_0500_),
    .B1(_1290_),
    .Y(_1291_));
 sky130_fd_sc_hd__a221oi_1 _4859_ (.A1(_0522_),
    .A2(_0492_),
    .B1(_0515_),
    .B2(_0496_),
    .C1(_1291_),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _4860_ (.A(_0514_),
    .B(_0486_),
    .Y(_1293_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(_0519_),
    .B(_0480_),
    .Y(_1294_));
 sky130_fd_sc_hd__or2_1 _4862_ (.A(_0896_),
    .B(_0525_),
    .X(_1295_));
 sky130_fd_sc_hd__o2111a_1 _4863_ (.A1(_1159_),
    .A2(_0511_),
    .B1(_1293_),
    .C1(_1294_),
    .D1(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__nand2_1 _4864_ (.A(_0538_),
    .B(_0707_),
    .Y(_1297_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(_0543_),
    .B(_0367_),
    .Y(_1298_));
 sky130_fd_sc_hd__nand2_1 _4866_ (.A(_1297_),
    .B(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__a221oi_1 _4867_ (.A1(_0377_),
    .A2(_0531_),
    .B1(_0709_),
    .B2(_0535_),
    .C1(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__and4_1 _4868_ (.A(_1289_),
    .B(_1292_),
    .C(_1296_),
    .D(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2_1 _4869_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1302_));
 sky130_fd_sc_hd__nand2_1 _4870_ (.A(_0562_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1303_));
 sky130_fd_sc_hd__or2_1 _4871_ (.A(_0605_),
    .B(_0567_),
    .X(_1304_));
 sky130_fd_sc_hd__o2111a_1 _4872_ (.A1(_0772_),
    .A2(_0554_),
    .B1(_1302_),
    .C1(_1303_),
    .D1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_0575_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1306_));
 sky130_fd_sc_hd__nand2_1 _4874_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1307_));
 sky130_fd_sc_hd__or2_1 _4875_ (.A(_0778_),
    .B(_0583_),
    .X(_1308_));
 sky130_fd_sc_hd__o2111a_1 _4876_ (.A1(_1058_),
    .A2(_0572_),
    .B1(_1306_),
    .C1(_1307_),
    .D1(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__or2_1 _4877_ (.A(_0767_),
    .B(_0596_),
    .X(_1310_));
 sky130_fd_sc_hd__o221a_1 _4878_ (.A1(_0565_),
    .A2(_0589_),
    .B1(_0764_),
    .B2(_0592_),
    .C1(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__o22ai_1 _4879_ (.A1(_1186_),
    .A2(_0607_),
    .B1(_0498_),
    .B2(_0610_),
    .Y(_1312_));
 sky130_fd_sc_hd__a221oi_1 _4880_ (.A1(_0504_),
    .A2(_0601_),
    .B1(_0520_),
    .B2(_0604_),
    .C1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__and4_1 _4881_ (.A(_1305_),
    .B(_1309_),
    .C(_1311_),
    .D(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__and3_1 _4882_ (.A(_1284_),
    .B(_1301_),
    .C(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__nand2_1 _4883_ (.A(_0618_),
    .B(_0549_),
    .Y(_1316_));
 sky130_fd_sc_hd__nand3_1 _4884_ (.A(_1253_),
    .B(_1315_),
    .C(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__inv_2 _4885_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_1318_));
 sky130_fd_sc_hd__a21oi_1 _4886_ (.A1(_1318_),
    .A2(_0932_),
    .B1(_2985_),
    .Y(_1319_));
 sky130_fd_sc_hd__o21a_1 _4887_ (.A1(_3103_),
    .A2(_1317_),
    .B1(_1319_),
    .X(_0292_));
 sky130_fd_sc_hd__inv_2 _4888_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1320_));
 sky130_fd_sc_hd__o22ai_1 _4889_ (.A1(_1195_),
    .A2(_3130_),
    .B1(_1320_),
    .B2(_3138_),
    .Y(_1321_));
 sky130_fd_sc_hd__a221oi_1 _4890_ (.A1(_0637_),
    .A2(_3115_),
    .B1(_0799_),
    .B2(_3122_),
    .C1(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_3160_),
    .B(_0632_),
    .Y(_1323_));
 sky130_fd_sc_hd__o21ai_1 _4892_ (.A1(_0634_),
    .A2(_3156_),
    .B1(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__a221oi_1 _4893_ (.A1(_0795_),
    .A2(_3147_),
    .B1(_3131_),
    .B2(_3152_),
    .C1(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(_3174_),
    .B(_3104_),
    .Y(_1326_));
 sky130_fd_sc_hd__nand2_1 _4895_ (.A(_3180_),
    .B(_3209_),
    .Y(_1327_));
 sky130_fd_sc_hd__or2_1 _4896_ (.A(_0787_),
    .B(_3187_),
    .X(_1328_));
 sky130_fd_sc_hd__o2111a_1 _4897_ (.A1(_1067_),
    .A2(_3169_),
    .B1(_1326_),
    .C1(_1327_),
    .D1(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_3202_),
    .B(_3301_),
    .Y(_1330_));
 sky130_fd_sc_hd__nand2_1 _4899_ (.A(_3208_),
    .B(_0661_),
    .Y(_1331_));
 sky130_fd_sc_hd__nand2_1 _4900_ (.A(_1330_),
    .B(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__a221oi_2 _4901_ (.A1(_0663_),
    .A2(_3194_),
    .B1(_0824_),
    .B2(_3198_),
    .C1(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__and4_1 _4902_ (.A(_1322_),
    .B(_1325_),
    .C(_1329_),
    .D(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__o22ai_1 _4903_ (.A1(_1210_),
    .A2(_3224_),
    .B1(_3236_),
    .B2(_3227_),
    .Y(_1335_));
 sky130_fd_sc_hd__a221oi_1 _4904_ (.A1(_3090_),
    .A2(_3218_),
    .B1(_3093_),
    .B2(_3221_),
    .C1(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_3241_),
    .B(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1337_));
 sky130_fd_sc_hd__o21ai_1 _4906_ (.A1(_0590_),
    .A2(_3238_),
    .B1(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__a221oi_1 _4907_ (.A1(_3096_),
    .A2(_3232_),
    .B1(_3099_),
    .B2(_3235_),
    .C1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__nand2_1 _4908_ (.A(_3256_),
    .B(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_1340_));
 sky130_fd_sc_hd__o21ai_1 _4909_ (.A1(_0643_),
    .A2(_3253_),
    .B1(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__a221oi_1 _4910_ (.A1(_3078_),
    .A2(_3247_),
    .B1(_3081_),
    .B2(_3250_),
    .C1(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__o22ai_1 _4911_ (.A1(_0587_),
    .A2(_3268_),
    .B1(_0594_),
    .B2(_3271_),
    .Y(_1343_));
 sky130_fd_sc_hd__a221oi_1 _4912_ (.A1(_0563_),
    .A2(_3262_),
    .B1(_0549_),
    .B2(_3265_),
    .C1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__and4_1 _4913_ (.A(_1336_),
    .B(_1339_),
    .C(_1342_),
    .D(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__o22ai_1 _4914_ (.A1(_0673_),
    .A2(_3288_),
    .B1(_0834_),
    .B2(_3291_),
    .Y(_1346_));
 sky130_fd_sc_hd__a221oi_1 _4915_ (.A1(_3366_),
    .A2(_3281_),
    .B1(_3370_),
    .B2(_3285_),
    .C1(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(_3296_),
    .B(_3323_),
    .Y(_1348_));
 sky130_fd_sc_hd__nand2_1 _4917_ (.A(_3300_),
    .B(_0831_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_1 _4918_ (.A(_3305_),
    .B(_0967_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4919_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1351_));
 sky130_fd_sc_hd__and4_1 _4920_ (.A(_1348_),
    .B(_1349_),
    .C(_1350_),
    .D(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__o22ai_1 _4921_ (.A1(_0658_),
    .A2(_3314_),
    .B1(_0820_),
    .B2(_3317_),
    .Y(_1353_));
 sky130_fd_sc_hd__a22o_1 _4922_ (.A1(_3320_),
    .A2(_0657_),
    .B1(_3322_),
    .B2(_0819_),
    .X(_1354_));
 sky130_fd_sc_hd__nor2_1 _4923_ (.A(_1353_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__inv_2 _4924_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .Y(_1356_));
 sky130_fd_sc_hd__o22ai_1 _4925_ (.A1(_1232_),
    .A2(_3336_),
    .B1(_1356_),
    .B2(_3339_),
    .Y(_1357_));
 sky130_fd_sc_hd__a221oi_1 _4926_ (.A1(_3391_),
    .A2(_3329_),
    .B1(_0686_),
    .B2(_3333_),
    .C1(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__and4_1 _4927_ (.A(_1347_),
    .B(_1352_),
    .C(_1355_),
    .D(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_3356_),
    .B(_0851_),
    .Y(_1360_));
 sky130_fd_sc_hd__nand2_1 _4929_ (.A(_3361_),
    .B(_0693_),
    .Y(_1361_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_1360_),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__a221oi_1 _4931_ (.A1(_3044_),
    .A2(_3349_),
    .B1(_3056_),
    .B2(_3353_),
    .C1(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_3375_),
    .B(_3357_),
    .Y(_1364_));
 sky130_fd_sc_hd__nand2_1 _4933_ (.A(_3380_),
    .B(_3362_),
    .Y(_1365_));
 sky130_fd_sc_hd__nand2_1 _4934_ (.A(_1364_),
    .B(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__a221oi_1 _4935_ (.A1(_3396_),
    .A2(_3369_),
    .B1(_0688_),
    .B2(_3372_),
    .C1(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__inv_2 _4936_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1368_));
 sky130_fd_sc_hd__nand2_1 _4937_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1369_));
 sky130_fd_sc_hd__nand2_1 _4938_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1370_));
 sky130_fd_sc_hd__or2_1 _4939_ (.A(_1117_),
    .B(_3400_),
    .X(_1371_));
 sky130_fd_sc_hd__o2111a_1 _4940_ (.A1(_1368_),
    .A2(_3387_),
    .B1(_1369_),
    .C1(_1370_),
    .D1(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__nand2_1 _4941_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_1373_));
 sky130_fd_sc_hd__o21ai_1 _4942_ (.A1(_3225_),
    .A2(_3413_),
    .B1(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__a221oi_1 _4943_ (.A1(_3059_),
    .A2(_3406_),
    .B1(_3062_),
    .B2(_3410_),
    .C1(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__and4_1 _4944_ (.A(_1363_),
    .B(_1367_),
    .C(_1372_),
    .D(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__and4_1 _4945_ (.A(_1334_),
    .B(_1345_),
    .C(_1359_),
    .D(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__nand2_1 _4946_ (.A(_0338_),
    .B(_0714_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _4947_ (.A(_0343_),
    .B(_0713_),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_1 _4948_ (.A(_1378_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__a221oi_1 _4949_ (.A1(_0869_),
    .A2(_0331_),
    .B1(_0448_),
    .B2(_0335_),
    .C1(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__inv_2 _4950_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_1382_));
 sky130_fd_sc_hd__o22ai_1 _4951_ (.A1(_1258_),
    .A2(_0350_),
    .B1(_1382_),
    .B2(_0353_),
    .Y(_1383_));
 sky130_fd_sc_hd__a22o_1 _4952_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .B1(_0359_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_1384_));
 sky130_fd_sc_hd__nor2_1 _4953_ (.A(_1383_),
    .B(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _4954_ (.A(_0376_),
    .B(_0339_),
    .Y(_1386_));
 sky130_fd_sc_hd__o21ai_1 _4955_ (.A1(_1001_),
    .A2(_0373_),
    .B1(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__a221oi_1 _4956_ (.A1(_0357_),
    .A2(_0366_),
    .B1(_0360_),
    .B2(_0370_),
    .C1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__nand2_1 _4957_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1389_));
 sky130_fd_sc_hd__o21ai_1 _4958_ (.A1(_0399_),
    .A2(_0391_),
    .B1(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__a221oi_1 _4959_ (.A1(_0434_),
    .A2(_0384_),
    .B1(_0438_),
    .B2(_0388_),
    .C1(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__and4_1 _4960_ (.A(_1381_),
    .B(_1385_),
    .C(_1388_),
    .D(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__nand2_1 _4961_ (.A(_0405_),
    .B(_0452_),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2_1 _4962_ (.A(_0409_),
    .B(_0427_),
    .Y(_1394_));
 sky130_fd_sc_hd__or2_1 _4963_ (.A(_0880_),
    .B(_0414_),
    .X(_1395_));
 sky130_fd_sc_hd__o2111a_1 _4964_ (.A1(_0417_),
    .A2(_0402_),
    .B1(_1393_),
    .C1(_1394_),
    .D1(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__nand2_1 _4965_ (.A(_0422_),
    .B(_0738_),
    .Y(_1397_));
 sky130_fd_sc_hd__nand2_1 _4966_ (.A(_0426_),
    .B(_0890_),
    .Y(_1398_));
 sky130_fd_sc_hd__or2_1 _4967_ (.A(_0460_),
    .B(_0431_),
    .X(_1399_));
 sky130_fd_sc_hd__o2111a_1 _4968_ (.A1(_0626_),
    .A2(_0419_),
    .B1(_1397_),
    .C1(_1398_),
    .D1(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_0447_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1401_));
 sky130_fd_sc_hd__o21ai_1 _4970_ (.A1(_0719_),
    .A2(_0444_),
    .B1(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__a221oi_1 _4971_ (.A1(_0874_),
    .A2(_0437_),
    .B1(_1012_),
    .B2(_0441_),
    .C1(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__nand2_1 _4972_ (.A(_0465_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1404_));
 sky130_fd_sc_hd__o21ai_1 _4973_ (.A1(_3183_),
    .A2(_0462_),
    .B1(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__a221oi_1 _4974_ (.A1(_3141_),
    .A2(_0455_),
    .B1(_3148_),
    .B2(_0459_),
    .C1(_1405_),
    .Y(_1406_));
 sky130_fd_sc_hd__and4_1 _4975_ (.A(_1396_),
    .B(_1400_),
    .C(_1403_),
    .D(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__and2_1 _4976_ (.A(_1392_),
    .B(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__inv_2 _4977_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .Y(_1409_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(_0479_),
    .B(_0532_),
    .Y(_1410_));
 sky130_fd_sc_hd__a22o_1 _4979_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_1411_));
 sky130_fd_sc_hd__inv_2 _4980_ (.A(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__o211a_1 _4981_ (.A1(_1409_),
    .A2(_0476_),
    .B1(_1410_),
    .C1(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__nand2_1 _4982_ (.A(_0503_),
    .B(_0480_),
    .Y(_1414_));
 sky130_fd_sc_hd__o21ai_1 _4983_ (.A1(_0472_),
    .A2(_0500_),
    .B1(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__a221oi_1 _4984_ (.A1(_0515_),
    .A2(_0492_),
    .B1(_0508_),
    .B2(_0496_),
    .C1(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__nand2_1 _4985_ (.A(_0514_),
    .B(_0544_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _4986_ (.A(_0519_),
    .B(_0745_),
    .Y(_1418_));
 sky130_fd_sc_hd__or2_1 _4987_ (.A(_1031_),
    .B(_0525_),
    .X(_1419_));
 sky130_fd_sc_hd__o2111a_1 _4988_ (.A1(_1285_),
    .A2(_0511_),
    .B1(_1417_),
    .C1(_1418_),
    .D1(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__nand2_1 _4989_ (.A(_0538_),
    .B(_0377_),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _4990_ (.A(_0543_),
    .B(_0707_),
    .Y(_1422_));
 sky130_fd_sc_hd__nand2_1 _4991_ (.A(_1421_),
    .B(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__a221oi_1 _4992_ (.A1(_0709_),
    .A2(_0531_),
    .B1(_0865_),
    .B2(_0535_),
    .C1(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__and4_1 _4993_ (.A(_1413_),
    .B(_1416_),
    .C(_1420_),
    .D(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__nand2_1 _4994_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1426_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_0562_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1427_));
 sky130_fd_sc_hd__or2_1 _4996_ (.A(_0608_),
    .B(_0567_),
    .X(_1428_));
 sky130_fd_sc_hd__o2111a_1 _4997_ (.A1(_0570_),
    .A2(_0554_),
    .B1(_1426_),
    .C1(_1427_),
    .D1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__nand2_1 _4998_ (.A(_0575_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_1 _4999_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1431_));
 sky130_fd_sc_hd__or2_1 _5000_ (.A(_0924_),
    .B(_0583_),
    .X(_1432_));
 sky130_fd_sc_hd__o2111a_1 _5001_ (.A1(_1186_),
    .A2(_0572_),
    .B1(_1430_),
    .C1(_1431_),
    .D1(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__or2_1 _5002_ (.A(_0581_),
    .B(_0596_),
    .X(_1434_));
 sky130_fd_sc_hd__o221a_1 _5003_ (.A1(_0767_),
    .A2(_0589_),
    .B1(_0565_),
    .B2(_0592_),
    .C1(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__o22ai_1 _5004_ (.A1(_0498_),
    .A2(_0607_),
    .B1(_0750_),
    .B2(_0610_),
    .Y(_1436_));
 sky130_fd_sc_hd__a221oi_1 _5005_ (.A1(_0520_),
    .A2(_0601_),
    .B1(_0522_),
    .B2(_0604_),
    .C1(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__and4_1 _5006_ (.A(_1429_),
    .B(_1433_),
    .C(_1435_),
    .D(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__and3_1 _5007_ (.A(_1408_),
    .B(_1425_),
    .C(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_0618_),
    .B(_0558_),
    .Y(_1440_));
 sky130_fd_sc_hd__nand3_1 _5009_ (.A(_1377_),
    .B(_1439_),
    .C(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__inv_2 _5010_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_1442_));
 sky130_fd_sc_hd__a21oi_1 _5011_ (.A1(_1442_),
    .A2(_0932_),
    .B1(_2985_),
    .Y(_1443_));
 sky130_fd_sc_hd__o21a_1 _5012_ (.A1(_3103_),
    .A2(_1441_),
    .B1(_1443_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _5013_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1444_));
 sky130_fd_sc_hd__o22ai_1 _5014_ (.A1(_1320_),
    .A2(_3130_),
    .B1(_1444_),
    .B2(_3138_),
    .Y(_1445_));
 sky130_fd_sc_hd__a221oi_1 _5015_ (.A1(_0799_),
    .A2(_3115_),
    .B1(_0661_),
    .B2(_3122_),
    .C1(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(_3160_),
    .B(_0795_),
    .Y(_1447_));
 sky130_fd_sc_hd__o21ai_1 _5017_ (.A1(_3165_),
    .A2(_3156_),
    .B1(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__a221oi_1 _5018_ (.A1(_3131_),
    .A2(_3147_),
    .B1(_3104_),
    .B2(_3152_),
    .C1(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__nand2_1 _5019_ (.A(_3174_),
    .B(_3116_),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _5020_ (.A(_3180_),
    .B(_3203_),
    .Y(_1451_));
 sky130_fd_sc_hd__or2_1 _5021_ (.A(_0934_),
    .B(_3187_),
    .X(_1452_));
 sky130_fd_sc_hd__o2111a_1 _5022_ (.A1(_1195_),
    .A2(_3169_),
    .B1(_1450_),
    .C1(_1451_),
    .D1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(_3202_),
    .B(_0663_),
    .Y(_1454_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(_3208_),
    .B(_3301_),
    .Y(_1455_));
 sky130_fd_sc_hd__nand2_1 _5025_ (.A(_1454_),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__a221oi_2 _5026_ (.A1(_0824_),
    .A2(_3194_),
    .B1(_0967_),
    .B2(_3198_),
    .C1(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__and4_1 _5027_ (.A(_1446_),
    .B(_1449_),
    .C(_1453_),
    .D(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__o22ai_1 _5028_ (.A1(_3236_),
    .A2(_3224_),
    .B1(_3266_),
    .B2(_3227_),
    .Y(_1459_));
 sky130_fd_sc_hd__a221oi_1 _5029_ (.A1(_3093_),
    .A2(_3218_),
    .B1(_3096_),
    .B2(_3221_),
    .C1(_1459_),
    .Y(_1460_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_3241_),
    .B(_0783_),
    .Y(_1461_));
 sky130_fd_sc_hd__o21ai_1 _5031_ (.A1(_0587_),
    .A2(_3238_),
    .B1(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__a221oi_1 _5032_ (.A1(_3099_),
    .A2(_3232_),
    .B1(_0619_),
    .B2(_3235_),
    .C1(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__nand2_1 _5033_ (.A(_3256_),
    .B(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1464_));
 sky130_fd_sc_hd__o21ai_1 _5034_ (.A1(_0805_),
    .A2(_3253_),
    .B1(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__a221oi_1 _5035_ (.A1(_3081_),
    .A2(_3247_),
    .B1(_3084_),
    .B2(_3250_),
    .C1(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__o22ai_1 _5036_ (.A1(_0594_),
    .A2(_3268_),
    .B1(_0775_),
    .B2(_3271_),
    .Y(_1467_));
 sky130_fd_sc_hd__a221oi_1 _5037_ (.A1(_0549_),
    .A2(_3262_),
    .B1(_0558_),
    .B2(_3265_),
    .C1(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__and4_1 _5038_ (.A(_1460_),
    .B(_1463_),
    .C(_1466_),
    .D(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__o22ai_1 _5039_ (.A1(_0834_),
    .A2(_3288_),
    .B1(_0975_),
    .B2(_3291_),
    .Y(_1470_));
 sky130_fd_sc_hd__a221oi_1 _5040_ (.A1(_3370_),
    .A2(_3281_),
    .B1(_3381_),
    .B2(_3285_),
    .C1(_1470_),
    .Y(_1471_));
 sky130_fd_sc_hd__nand2_1 _5041_ (.A(_3296_),
    .B(_0670_),
    .Y(_1472_));
 sky130_fd_sc_hd__nand2_1 _5042_ (.A(_3300_),
    .B(_3275_),
    .Y(_1473_));
 sky130_fd_sc_hd__nand2_1 _5043_ (.A(_3305_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _5044_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_1475_));
 sky130_fd_sc_hd__and4_1 _5045_ (.A(_1472_),
    .B(_1473_),
    .C(_1474_),
    .D(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__o22ai_1 _5046_ (.A1(_0820_),
    .A2(_3314_),
    .B1(_3334_),
    .B2(_3317_),
    .Y(_1477_));
 sky130_fd_sc_hd__a22o_1 _5047_ (.A1(_3320_),
    .A2(_0819_),
    .B1(_3322_),
    .B2(_3326_),
    .X(_1478_));
 sky130_fd_sc_hd__nor2_1 _5048_ (.A(_1477_),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__inv_2 _5049_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_1480_));
 sky130_fd_sc_hd__o22ai_1 _5050_ (.A1(_1356_),
    .A2(_3336_),
    .B1(_1480_),
    .B2(_3339_),
    .Y(_1481_));
 sky130_fd_sc_hd__a221oi_1 _5051_ (.A1(_0686_),
    .A2(_3329_),
    .B1(_3396_),
    .B2(_3333_),
    .C1(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__and4_1 _5052_ (.A(_1471_),
    .B(_1476_),
    .C(_1479_),
    .D(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_1 _5053_ (.A(_3356_),
    .B(_3044_),
    .Y(_1484_));
 sky130_fd_sc_hd__nand2_1 _5054_ (.A(_3361_),
    .B(_0851_),
    .Y(_1485_));
 sky130_fd_sc_hd__nand2_1 _5055_ (.A(_1484_),
    .B(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__a221oi_1 _5056_ (.A1(_3056_),
    .A2(_3349_),
    .B1(_3059_),
    .B2(_3353_),
    .C1(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__nand2_1 _5057_ (.A(_3375_),
    .B(_3343_),
    .Y(_1488_));
 sky130_fd_sc_hd__nand2_1 _5058_ (.A(_3380_),
    .B(_3357_),
    .Y(_1489_));
 sky130_fd_sc_hd__nand2_1 _5059_ (.A(_1488_),
    .B(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__a221oi_1 _5060_ (.A1(_0688_),
    .A2(_3369_),
    .B1(_3362_),
    .B2(_3372_),
    .C1(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__inv_2 _5061_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_1 _5062_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1493_));
 sky130_fd_sc_hd__nand2_1 _5063_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1494_));
 sky130_fd_sc_hd__or2_1 _5064_ (.A(_1244_),
    .B(_3400_),
    .X(_1495_));
 sky130_fd_sc_hd__o2111a_1 _5065_ (.A1(_1492_),
    .A2(_3387_),
    .B1(_1493_),
    .C1(_1494_),
    .D1(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__nand2_1 _5066_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_1497_));
 sky130_fd_sc_hd__o21ai_1 _5067_ (.A1(_0643_),
    .A2(_3413_),
    .B1(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__a221oi_1 _5068_ (.A1(_3062_),
    .A2(_3406_),
    .B1(_3065_),
    .B2(_3410_),
    .C1(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__and4_1 _5069_ (.A(_1487_),
    .B(_1491_),
    .C(_1496_),
    .D(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__and4_1 _5070_ (.A(_1458_),
    .B(_1469_),
    .C(_1483_),
    .D(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_0338_),
    .B(_0869_),
    .Y(_1502_));
 sky130_fd_sc_hd__nand2_1 _5072_ (.A(_0343_),
    .B(_0714_),
    .Y(_1503_));
 sky130_fd_sc_hd__nand2_1 _5073_ (.A(_1502_),
    .B(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__a221oi_1 _5074_ (.A1(_0448_),
    .A2(_0331_),
    .B1(_0434_),
    .B2(_0335_),
    .C1(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__inv_2 _5075_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1506_));
 sky130_fd_sc_hd__o22ai_1 _5076_ (.A1(_1382_),
    .A2(_0350_),
    .B1(_1506_),
    .B2(_0353_),
    .Y(_1507_));
 sky130_fd_sc_hd__a22o_1 _5077_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .B1(_0359_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_1508_));
 sky130_fd_sc_hd__nor2_1 _5078_ (.A(_1507_),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _5079_ (.A(_0376_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1510_));
 sky130_fd_sc_hd__o21ai_1 _5080_ (.A1(_1131_),
    .A2(_0373_),
    .B1(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__a221oi_1 _5081_ (.A1(_0360_),
    .A2(_0366_),
    .B1(_0344_),
    .B2(_0370_),
    .C1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1513_));
 sky130_fd_sc_hd__o21ai_1 _5083_ (.A1(_0719_),
    .A2(_0391_),
    .B1(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__a221oi_1 _5084_ (.A1(_0438_),
    .A2(_0384_),
    .B1(_0410_),
    .B2(_0388_),
    .C1(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__and4_1 _5085_ (.A(_1505_),
    .B(_1509_),
    .C(_1512_),
    .D(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_0405_),
    .B(_0456_),
    .Y(_1517_));
 sky130_fd_sc_hd__nand2_1 _5087_ (.A(_0409_),
    .B(_0729_),
    .Y(_1518_));
 sky130_fd_sc_hd__or2_1 _5088_ (.A(_1017_),
    .B(_0414_),
    .X(_1519_));
 sky130_fd_sc_hd__o2111a_1 _5089_ (.A1(_0727_),
    .A2(_0402_),
    .B1(_1517_),
    .C1(_1518_),
    .D1(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__nand2_1 _5090_ (.A(_0422_),
    .B(_0889_),
    .Y(_1521_));
 sky130_fd_sc_hd__nand2_1 _5091_ (.A(_0426_),
    .B(_3161_),
    .Y(_1522_));
 sky130_fd_sc_hd__or2_1 _5092_ (.A(_3153_),
    .B(_0431_),
    .X(_1523_));
 sky130_fd_sc_hd__o2111a_1 _5093_ (.A1(_0790_),
    .A2(_0419_),
    .B1(_1521_),
    .C1(_1522_),
    .D1(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_0447_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1525_));
 sky130_fd_sc_hd__o21ai_1 _5095_ (.A1(_0412_),
    .A2(_0444_),
    .B1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__a221oi_1 _5096_ (.A1(_1012_),
    .A2(_0437_),
    .B1(_0427_),
    .B2(_0441_),
    .C1(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__nand2_1 _5097_ (.A(_0465_),
    .B(_0630_),
    .Y(_1528_));
 sky130_fd_sc_hd__o21ai_1 _5098_ (.A1(_0634_),
    .A2(_0462_),
    .B1(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__a221oi_1 _5099_ (.A1(_3148_),
    .A2(_0455_),
    .B1(_3175_),
    .B2(_0459_),
    .C1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__and4_1 _5100_ (.A(_1520_),
    .B(_1524_),
    .C(_1527_),
    .D(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__and2_1 _5101_ (.A(_1516_),
    .B(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__inv_2 _5102_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .Y(_1533_));
 sky130_fd_sc_hd__nand2_1 _5103_ (.A(_0479_),
    .B(_0363_),
    .Y(_1534_));
 sky130_fd_sc_hd__a22o_1 _5104_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_1535_));
 sky130_fd_sc_hd__inv_2 _5105_ (.A(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__o211a_1 _5106_ (.A1(_1533_),
    .A2(_0476_),
    .B1(_1534_),
    .C1(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__nand2_1 _5107_ (.A(_0503_),
    .B(_0745_),
    .Y(_1538_));
 sky130_fd_sc_hd__o21ai_1 _5108_ (.A1(_0744_),
    .A2(_0500_),
    .B1(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__a221oi_1 _5109_ (.A1(_0508_),
    .A2(_0492_),
    .B1(_0471_),
    .B2(_0496_),
    .C1(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__nand2_1 _5110_ (.A(_0514_),
    .B(_0539_),
    .Y(_1541_));
 sky130_fd_sc_hd__nand2_1 _5111_ (.A(_0519_),
    .B(_0486_),
    .Y(_1542_));
 sky130_fd_sc_hd__or2_1 _5112_ (.A(_1159_),
    .B(_0525_),
    .X(_1543_));
 sky130_fd_sc_hd__o2111a_1 _5113_ (.A1(_1409_),
    .A2(_0511_),
    .B1(_1541_),
    .C1(_1542_),
    .D1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__nand2_1 _5114_ (.A(_0538_),
    .B(_0709_),
    .Y(_1545_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_0543_),
    .B(_0377_),
    .Y(_1546_));
 sky130_fd_sc_hd__nand2_1 _5116_ (.A(_1545_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__a221oi_1 _5117_ (.A1(_0865_),
    .A2(_0531_),
    .B1(_0357_),
    .B2(_0535_),
    .C1(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__and4_1 _5118_ (.A(_1537_),
    .B(_1540_),
    .C(_1544_),
    .D(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__nand2_1 _5119_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1550_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_0562_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1551_));
 sky130_fd_sc_hd__or2_1 _5121_ (.A(_0778_),
    .B(_0567_),
    .X(_1552_));
 sky130_fd_sc_hd__o2111a_1 _5122_ (.A1(_0605_),
    .A2(_0554_),
    .B1(_1550_),
    .C1(_1551_),
    .D1(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__nand2_1 _5123_ (.A(_0575_),
    .B(_0493_),
    .Y(_1554_));
 sky130_fd_sc_hd__nand2_1 _5124_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1555_));
 sky130_fd_sc_hd__or2_1 _5125_ (.A(_1058_),
    .B(_0583_),
    .X(_1556_));
 sky130_fd_sc_hd__o2111a_1 _5126_ (.A1(_0498_),
    .A2(_0572_),
    .B1(_1554_),
    .C1(_1555_),
    .D1(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__or2_1 _5127_ (.A(_0772_),
    .B(_0596_),
    .X(_1558_));
 sky130_fd_sc_hd__o221a_1 _5128_ (.A1(_0581_),
    .A2(_0589_),
    .B1(_0767_),
    .B2(_0592_),
    .C1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__o22ai_1 _5129_ (.A1(_0750_),
    .A2(_0607_),
    .B1(_0901_),
    .B2(_0610_),
    .Y(_1560_));
 sky130_fd_sc_hd__a221oi_1 _5130_ (.A1(_0522_),
    .A2(_0601_),
    .B1(_0515_),
    .B2(_0604_),
    .C1(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__and4_1 _5131_ (.A(_1553_),
    .B(_1557_),
    .C(_1559_),
    .D(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__and3_1 _5132_ (.A(_1532_),
    .B(_1549_),
    .C(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(_0618_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_1564_));
 sky130_fd_sc_hd__nand3_1 _5134_ (.A(_1501_),
    .B(_1563_),
    .C(_1564_),
    .Y(_1565_));
 sky130_fd_sc_hd__inv_2 _5135_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_1566_));
 sky130_fd_sc_hd__a21oi_1 _5136_ (.A1(_1566_),
    .A2(_3102_),
    .B1(_2985_),
    .Y(_1567_));
 sky130_fd_sc_hd__o21a_1 _5137_ (.A1(_3103_),
    .A2(_1565_),
    .B1(_1567_),
    .X(_0290_));
 sky130_fd_sc_hd__inv_2 _5138_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1568_));
 sky130_fd_sc_hd__o22ai_1 _5139_ (.A1(_1444_),
    .A2(_3130_),
    .B1(_1568_),
    .B2(_3138_),
    .Y(_1569_));
 sky130_fd_sc_hd__a221oi_1 _5140_ (.A1(_0661_),
    .A2(_3115_),
    .B1(_3301_),
    .B2(_3122_),
    .C1(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__nand2_1 _5141_ (.A(_3160_),
    .B(_3131_),
    .Y(_1571_));
 sky130_fd_sc_hd__o21ai_1 _5142_ (.A1(_3123_),
    .A2(_3156_),
    .B1(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__a221oi_1 _5143_ (.A1(_3104_),
    .A2(_3147_),
    .B1(_3116_),
    .B2(_3152_),
    .C1(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2_1 _5144_ (.A(_3174_),
    .B(_3209_),
    .Y(_1574_));
 sky130_fd_sc_hd__nand2_1 _5145_ (.A(_3180_),
    .B(_3190_),
    .Y(_1575_));
 sky130_fd_sc_hd__or2_1 _5146_ (.A(_1067_),
    .B(_3187_),
    .X(_1576_));
 sky130_fd_sc_hd__o2111a_1 _5147_ (.A1(_1320_),
    .A2(_3169_),
    .B1(_1574_),
    .C1(_1575_),
    .D1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__nand2_1 _5148_ (.A(_3202_),
    .B(_0824_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_3208_),
    .B(_0663_),
    .Y(_1579_));
 sky130_fd_sc_hd__nand2_1 _5150_ (.A(_1578_),
    .B(_1579_),
    .Y(_1580_));
 sky130_fd_sc_hd__a221oi_1 _5151_ (.A1(_0967_),
    .A2(_3194_),
    .B1(_3323_),
    .B2(_3198_),
    .C1(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__and4_1 _5152_ (.A(_1570_),
    .B(_1573_),
    .C(_1577_),
    .D(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__o22ai_1 _5153_ (.A1(_3266_),
    .A2(_3224_),
    .B1(_3269_),
    .B2(_3227_),
    .Y(_1583_));
 sky130_fd_sc_hd__a221oi_1 _5154_ (.A1(_3096_),
    .A2(_3218_),
    .B1(_3099_),
    .B2(_3221_),
    .C1(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_3241_),
    .B(_0586_),
    .Y(_1585_));
 sky130_fd_sc_hd__o21ai_1 _5156_ (.A1(_0594_),
    .A2(_3238_),
    .B1(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__a221oi_1 _5157_ (.A1(_0619_),
    .A2(_3232_),
    .B1(_0783_),
    .B2(_3235_),
    .C1(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__nand2_1 _5158_ (.A(_3256_),
    .B(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1588_));
 sky130_fd_sc_hd__o21ai_1 _5159_ (.A1(_0950_),
    .A2(_3253_),
    .B1(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__a221oi_1 _5160_ (.A1(_3084_),
    .A2(_3247_),
    .B1(_3087_),
    .B2(_3250_),
    .C1(_1589_),
    .Y(_1590_));
 sky130_fd_sc_hd__o22ai_1 _5161_ (.A1(_0775_),
    .A2(_3268_),
    .B1(_0550_),
    .B2(_3271_),
    .Y(_1591_));
 sky130_fd_sc_hd__a221oi_1 _5162_ (.A1(_0558_),
    .A2(_3262_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .B2(_3265_),
    .C1(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__and4_1 _5163_ (.A(_1584_),
    .B(_1587_),
    .C(_1590_),
    .D(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__o22ai_1 _5164_ (.A1(_0975_),
    .A2(_3288_),
    .B1(_1105_),
    .B2(_3291_),
    .Y(_1594_));
 sky130_fd_sc_hd__a221oi_1 _5165_ (.A1(_3381_),
    .A2(_3281_),
    .B1(_3376_),
    .B2(_3285_),
    .C1(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__nand2_1 _5166_ (.A(_3296_),
    .B(_0831_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _5167_ (.A(_3300_),
    .B(_3282_),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _5168_ (.A(_3305_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_1 _5169_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_1599_));
 sky130_fd_sc_hd__and4_1 _5170_ (.A(_1596_),
    .B(_1597_),
    .C(_1598_),
    .D(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__o22ai_1 _5171_ (.A1(_3334_),
    .A2(_3314_),
    .B1(_3337_),
    .B2(_3317_),
    .Y(_1601_));
 sky130_fd_sc_hd__a22o_1 _5172_ (.A1(_3320_),
    .A2(_3326_),
    .B1(_3322_),
    .B2(_3330_),
    .X(_1602_));
 sky130_fd_sc_hd__nor2_1 _5173_ (.A(_1601_),
    .B(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__o22ai_1 _5174_ (.A1(_1480_),
    .A2(_3336_),
    .B1(_3398_),
    .B2(_3339_),
    .Y(_1604_));
 sky130_fd_sc_hd__a221oi_1 _5175_ (.A1(_3396_),
    .A2(_3329_),
    .B1(_0688_),
    .B2(_3333_),
    .C1(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__and4_1 _5176_ (.A(_1595_),
    .B(_1600_),
    .C(_1603_),
    .D(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__nand2_1 _5177_ (.A(_3356_),
    .B(_3056_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(_3361_),
    .B(_3044_),
    .Y(_1608_));
 sky130_fd_sc_hd__nand2_1 _5179_ (.A(_1607_),
    .B(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__a221oi_1 _5180_ (.A1(_3059_),
    .A2(_3349_),
    .B1(_3062_),
    .B2(_3353_),
    .C1(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__nand2_1 _5181_ (.A(_3375_),
    .B(_3350_),
    .Y(_1611_));
 sky130_fd_sc_hd__nand2_1 _5182_ (.A(_3380_),
    .B(_3343_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _5183_ (.A(_1611_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__a221oi_1 _5184_ (.A1(_3362_),
    .A2(_3369_),
    .B1(_3357_),
    .B2(_3372_),
    .C1(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__nand2_1 _5185_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2_1 _5186_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1616_));
 sky130_fd_sc_hd__or2_1 _5187_ (.A(_1368_),
    .B(_3400_),
    .X(_1617_));
 sky130_fd_sc_hd__o2111a_1 _5188_ (.A1(_3411_),
    .A2(_3387_),
    .B1(_1615_),
    .C1(_1616_),
    .D1(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1619_));
 sky130_fd_sc_hd__o21ai_1 _5190_ (.A1(_0805_),
    .A2(_3413_),
    .B1(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__a221oi_1 _5191_ (.A1(_3065_),
    .A2(_3406_),
    .B1(_3068_),
    .B2(_3410_),
    .C1(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__and4_1 _5192_ (.A(_1610_),
    .B(_1614_),
    .C(_1618_),
    .D(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__and4_1 _5193_ (.A(_1582_),
    .B(_1593_),
    .C(_1606_),
    .D(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__nand2_1 _5194_ (.A(_0338_),
    .B(_0448_),
    .Y(_1624_));
 sky130_fd_sc_hd__nand2_1 _5195_ (.A(_0343_),
    .B(_0869_),
    .Y(_1625_));
 sky130_fd_sc_hd__nand2_1 _5196_ (.A(_1624_),
    .B(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__a221oi_1 _5197_ (.A1(_0434_),
    .A2(_0331_),
    .B1(_0438_),
    .B2(_0335_),
    .C1(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__inv_2 _5198_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1628_));
 sky130_fd_sc_hd__o22ai_1 _5199_ (.A1(_1506_),
    .A2(_0350_),
    .B1(_1628_),
    .B2(_0353_),
    .Y(_1629_));
 sky130_fd_sc_hd__a22o_1 _5200_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .B1(_0359_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_1630_));
 sky130_fd_sc_hd__nor2_1 _5201_ (.A(_1629_),
    .B(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__nand2_1 _5202_ (.A(_0376_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_1632_));
 sky130_fd_sc_hd__o21ai_1 _5203_ (.A1(_1258_),
    .A2(_0373_),
    .B1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__a221oi_1 _5204_ (.A1(_0344_),
    .A2(_0366_),
    .B1(_0339_),
    .B2(_0370_),
    .C1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__nand2_1 _5205_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1635_));
 sky130_fd_sc_hd__o21ai_1 _5206_ (.A1(_0412_),
    .A2(_0391_),
    .B1(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__a221oi_1 _5207_ (.A1(_0410_),
    .A2(_0384_),
    .B1(_0722_),
    .B2(_0388_),
    .C1(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__and4_1 _5208_ (.A(_1627_),
    .B(_1631_),
    .C(_1634_),
    .D(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__nand2_1 _5209_ (.A(_0405_),
    .B(_0738_),
    .Y(_1639_));
 sky130_fd_sc_hd__nand2_1 _5210_ (.A(_0409_),
    .B(_0452_),
    .Y(_1640_));
 sky130_fd_sc_hd__or2_1 _5211_ (.A(_0460_),
    .B(_0414_),
    .X(_1641_));
 sky130_fd_sc_hd__o2111a_1 _5212_ (.A1(_0880_),
    .A2(_0402_),
    .B1(_1639_),
    .C1(_1640_),
    .D1(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__nand2_1 _5213_ (.A(_0422_),
    .B(_0890_),
    .Y(_1643_));
 sky130_fd_sc_hd__nand2_1 _5214_ (.A(_0426_),
    .B(_3141_),
    .Y(_1644_));
 sky130_fd_sc_hd__or2_1 _5215_ (.A(_0626_),
    .B(_0431_),
    .X(_1645_));
 sky130_fd_sc_hd__o2111a_1 _5216_ (.A1(_0937_),
    .A2(_0419_),
    .B1(_1643_),
    .C1(_1644_),
    .D1(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_1 _5217_ (.A(_0447_),
    .B(_1012_),
    .Y(_1647_));
 sky130_fd_sc_hd__o21ai_1 _5218_ (.A1(_0724_),
    .A2(_0444_),
    .B1(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__a221oi_1 _5219_ (.A1(_0427_),
    .A2(_0437_),
    .B1(_0729_),
    .B2(_0441_),
    .C1(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(_0465_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1650_));
 sky130_fd_sc_hd__o21ai_1 _5221_ (.A1(_3165_),
    .A2(_0462_),
    .B1(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__a221oi_1 _5222_ (.A1(_3175_),
    .A2(_0455_),
    .B1(_0630_),
    .B2(_0459_),
    .C1(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__and4_1 _5223_ (.A(_1642_),
    .B(_1646_),
    .C(_1649_),
    .D(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__and2_1 _5224_ (.A(_1638_),
    .B(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__inv_2 _5225_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_1655_));
 sky130_fd_sc_hd__nand2_1 _5226_ (.A(_0479_),
    .B(_0367_),
    .Y(_1656_));
 sky130_fd_sc_hd__a22o_1 _5227_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_1657_));
 sky130_fd_sc_hd__inv_2 _5228_ (.A(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__o211a_1 _5229_ (.A1(_1655_),
    .A2(_0476_),
    .B1(_1656_),
    .C1(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__nand2_1 _5230_ (.A(_0503_),
    .B(_0486_),
    .Y(_1660_));
 sky130_fd_sc_hd__o21ai_1 _5231_ (.A1(_0896_),
    .A2(_0500_),
    .B1(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__a221oi_1 _5232_ (.A1(_0471_),
    .A2(_0492_),
    .B1(_0480_),
    .B2(_0496_),
    .C1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_0514_),
    .B(_0528_),
    .Y(_1663_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(_0519_),
    .B(_0544_),
    .Y(_1664_));
 sky130_fd_sc_hd__or2_1 _5235_ (.A(_1285_),
    .B(_0525_),
    .X(_1665_));
 sky130_fd_sc_hd__o2111a_1 _5236_ (.A1(_1533_),
    .A2(_0511_),
    .B1(_1663_),
    .C1(_1664_),
    .D1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__nand2_1 _5237_ (.A(_0538_),
    .B(_0865_),
    .Y(_1667_));
 sky130_fd_sc_hd__nand2_1 _5238_ (.A(_0543_),
    .B(_0709_),
    .Y(_1668_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(_1667_),
    .B(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__a221oi_1 _5240_ (.A1(_0357_),
    .A2(_0531_),
    .B1(_0360_),
    .B2(_0535_),
    .C1(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__and4_1 _5241_ (.A(_1659_),
    .B(_1662_),
    .C(_1666_),
    .D(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1672_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_0562_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1673_));
 sky130_fd_sc_hd__or2_1 _5244_ (.A(_0924_),
    .B(_0567_),
    .X(_1674_));
 sky130_fd_sc_hd__o2111a_1 _5245_ (.A1(_0608_),
    .A2(_0554_),
    .B1(_1672_),
    .C1(_1673_),
    .D1(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__nand2_1 _5246_ (.A(_0575_),
    .B(_0497_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1677_));
 sky130_fd_sc_hd__or2_1 _5248_ (.A(_1186_),
    .B(_0583_),
    .X(_1678_));
 sky130_fd_sc_hd__o2111a_1 _5249_ (.A1(_0750_),
    .A2(_0572_),
    .B1(_1676_),
    .C1(_1677_),
    .D1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(_0570_),
    .B(_0596_),
    .X(_1680_));
 sky130_fd_sc_hd__o221a_1 _5251_ (.A1(_0772_),
    .A2(_0589_),
    .B1(_0581_),
    .B2(_0592_),
    .C1(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__o22ai_1 _5252_ (.A1(_0901_),
    .A2(_0607_),
    .B1(_0523_),
    .B2(_0610_),
    .Y(_1682_));
 sky130_fd_sc_hd__a221oi_1 _5253_ (.A1(_0515_),
    .A2(_0601_),
    .B1(_0508_),
    .B2(_0604_),
    .C1(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__and4_1 _5254_ (.A(_1675_),
    .B(_1679_),
    .C(_1681_),
    .D(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__and3_1 _5255_ (.A(_1654_),
    .B(_1671_),
    .C(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(_0618_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_1686_));
 sky130_fd_sc_hd__nand3_1 _5257_ (.A(_1623_),
    .B(_1685_),
    .C(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__inv_2 _5258_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_1688_));
 sky130_fd_sc_hd__a21oi_1 _5259_ (.A1(_1688_),
    .A2(_3102_),
    .B1(_2985_),
    .Y(_1689_));
 sky130_fd_sc_hd__o21a_1 _5260_ (.A1(_3103_),
    .A2(_1687_),
    .B1(_1689_),
    .X(_0289_));
 sky130_fd_sc_hd__inv_2 _5261_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1690_));
 sky130_fd_sc_hd__o22ai_1 _5262_ (.A1(_1568_),
    .A2(_3130_),
    .B1(_1690_),
    .B2(_3138_),
    .Y(_1691_));
 sky130_fd_sc_hd__a221oi_1 _5263_ (.A1(_3301_),
    .A2(_3115_),
    .B1(_0663_),
    .B2(_3122_),
    .C1(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__nand2_1 _5264_ (.A(_3160_),
    .B(_3104_),
    .Y(_1693_));
 sky130_fd_sc_hd__o21ai_1 _5265_ (.A1(_3132_),
    .A2(_3156_),
    .B1(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__a221oi_2 _5266_ (.A1(_3116_),
    .A2(_3147_),
    .B1(_3209_),
    .B2(_3152_),
    .C1(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand2_1 _5267_ (.A(_3174_),
    .B(_3203_),
    .Y(_1696_));
 sky130_fd_sc_hd__nand2_1 _5268_ (.A(_3180_),
    .B(_3195_),
    .Y(_1697_));
 sky130_fd_sc_hd__or2_1 _5269_ (.A(_1195_),
    .B(_3187_),
    .X(_1698_));
 sky130_fd_sc_hd__o2111a_1 _5270_ (.A1(_1444_),
    .A2(_3169_),
    .B1(_1696_),
    .C1(_1697_),
    .D1(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__nand2_1 _5271_ (.A(_3202_),
    .B(_0967_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand2_1 _5272_ (.A(_3208_),
    .B(_0824_),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _5273_ (.A(_1700_),
    .B(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__a221oi_1 _5274_ (.A1(_3323_),
    .A2(_3194_),
    .B1(_0670_),
    .B2(_3198_),
    .C1(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__and4_1 _5275_ (.A(_1692_),
    .B(_1695_),
    .C(_1699_),
    .D(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__o22ai_1 _5276_ (.A1(_3269_),
    .A2(_3224_),
    .B1(_0653_),
    .B2(_3227_),
    .Y(_1705_));
 sky130_fd_sc_hd__a221oi_1 _5277_ (.A1(_3099_),
    .A2(_3218_),
    .B1(_0619_),
    .B2(_3221_),
    .C1(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__nand2_1 _5278_ (.A(_3241_),
    .B(_0593_),
    .Y(_1707_));
 sky130_fd_sc_hd__o21ai_1 _5279_ (.A1(_0775_),
    .A2(_3238_),
    .B1(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__a221oi_1 _5280_ (.A1(_0783_),
    .A2(_3232_),
    .B1(_0586_),
    .B2(_3235_),
    .C1(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_1 _5281_ (.A(_3256_),
    .B(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1710_));
 sky130_fd_sc_hd__o21ai_1 _5282_ (.A1(_1083_),
    .A2(_3253_),
    .B1(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__a221oi_1 _5283_ (.A1(_3087_),
    .A2(_3247_),
    .B1(_3090_),
    .B2(_3250_),
    .C1(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__o22ai_1 _5284_ (.A1(_0550_),
    .A2(_3268_),
    .B1(_0764_),
    .B2(_3271_),
    .Y(_1713_));
 sky130_fd_sc_hd__a221oi_1 _5285_ (.A1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .A2(_3262_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .B2(_3265_),
    .C1(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__and4_1 _5286_ (.A(_1706_),
    .B(_1709_),
    .C(_1712_),
    .D(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__o22ai_1 _5287_ (.A1(_1105_),
    .A2(_3288_),
    .B1(_1232_),
    .B2(_3291_),
    .Y(_1716_));
 sky130_fd_sc_hd__a221oi_1 _5288_ (.A1(_3376_),
    .A2(_3281_),
    .B1(_3391_),
    .B2(_3285_),
    .C1(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hd__nand2_1 _5289_ (.A(_3296_),
    .B(_3275_),
    .Y(_1718_));
 sky130_fd_sc_hd__nand2_1 _5290_ (.A(_3300_),
    .B(_0657_),
    .Y(_1719_));
 sky130_fd_sc_hd__nand2_1 _5291_ (.A(_3305_),
    .B(_0831_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand2_1 _5292_ (.A(_3309_),
    .B(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_1721_));
 sky130_fd_sc_hd__and4_1 _5293_ (.A(_1718_),
    .B(_1719_),
    .C(_1720_),
    .D(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__o22ai_1 _5294_ (.A1(_3337_),
    .A2(_3314_),
    .B1(_0673_),
    .B2(_3317_),
    .Y(_1723_));
 sky130_fd_sc_hd__a22o_1 _5295_ (.A1(_3320_),
    .A2(_3330_),
    .B1(_3322_),
    .B2(_3366_),
    .X(_1724_));
 sky130_fd_sc_hd__nor2_1 _5296_ (.A(_1723_),
    .B(_1724_),
    .Y(_1725_));
 sky130_fd_sc_hd__o22ai_1 _5297_ (.A1(_3398_),
    .A2(_3336_),
    .B1(_0690_),
    .B2(_3339_),
    .Y(_1726_));
 sky130_fd_sc_hd__a221oi_1 _5298_ (.A1(_0688_),
    .A2(_3329_),
    .B1(_3362_),
    .B2(_3333_),
    .C1(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__and4_1 _5299_ (.A(_1717_),
    .B(_1722_),
    .C(_1725_),
    .D(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(_3356_),
    .B(_3059_),
    .Y(_1729_));
 sky130_fd_sc_hd__nand2_1 _5301_ (.A(_3361_),
    .B(_3056_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_1 _5302_ (.A(_1729_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__a221oi_1 _5303_ (.A1(_3062_),
    .A2(_3349_),
    .B1(_3065_),
    .B2(_3353_),
    .C1(_1731_),
    .Y(_1732_));
 sky130_fd_sc_hd__nand2_1 _5304_ (.A(_3375_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _5305_ (.A(_3380_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(_1733_),
    .B(_1734_),
    .Y(_1735_));
 sky130_fd_sc_hd__a221oi_1 _5307_ (.A1(_3357_),
    .A2(_3369_),
    .B1(_3343_),
    .B2(_3372_),
    .C1(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2_1 _5308_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1737_));
 sky130_fd_sc_hd__nand2_1 _5309_ (.A(_3395_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_1738_));
 sky130_fd_sc_hd__or2_1 _5310_ (.A(_1492_),
    .B(_3400_),
    .X(_1739_));
 sky130_fd_sc_hd__o2111a_1 _5311_ (.A1(_3251_),
    .A2(_3387_),
    .B1(_1737_),
    .C1(_1738_),
    .D1(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__nand2_1 _5312_ (.A(_3416_),
    .B(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_1741_));
 sky130_fd_sc_hd__o21ai_1 _5313_ (.A1(_0950_),
    .A2(_3413_),
    .B1(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__a221oi_1 _5314_ (.A1(_3068_),
    .A2(_3406_),
    .B1(_3071_),
    .B2(_3410_),
    .C1(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hd__and4_1 _5315_ (.A(_1732_),
    .B(_1736_),
    .C(_1740_),
    .D(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__and4_1 _5316_ (.A(_1704_),
    .B(_1715_),
    .C(_1728_),
    .D(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__nand2_1 _5317_ (.A(_0338_),
    .B(_0434_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5318_ (.A(_0343_),
    .B(_0448_),
    .Y(_1747_));
 sky130_fd_sc_hd__nand2_1 _5319_ (.A(_1746_),
    .B(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__a221oi_1 _5320_ (.A1(_0438_),
    .A2(_0331_),
    .B1(_0410_),
    .B2(_0335_),
    .C1(_1748_),
    .Y(_1749_));
 sky130_fd_sc_hd__inv_2 _5321_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1750_));
 sky130_fd_sc_hd__o22ai_1 _5322_ (.A1(_1628_),
    .A2(_0350_),
    .B1(_1750_),
    .B2(_0353_),
    .Y(_1751_));
 sky130_fd_sc_hd__a22o_1 _5323_ (.A1(_0356_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .B1(_0359_),
    .B2(_0869_),
    .X(_1752_));
 sky130_fd_sc_hd__nor2_1 _5324_ (.A(_1751_),
    .B(_1752_),
    .Y(_1753_));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(_0376_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1754_));
 sky130_fd_sc_hd__o21ai_1 _5326_ (.A1(_1382_),
    .A2(_0373_),
    .B1(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__a221oi_2 _5327_ (.A1(_0339_),
    .A2(_0366_),
    .B1(_0326_),
    .B2(_0370_),
    .C1(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _5328_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1757_));
 sky130_fd_sc_hd__o21ai_1 _5329_ (.A1(_0724_),
    .A2(_0391_),
    .B1(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__a221oi_1 _5330_ (.A1(_0722_),
    .A2(_0384_),
    .B1(_0876_),
    .B2(_0388_),
    .C1(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__and4_1 _5331_ (.A(_1749_),
    .B(_1753_),
    .C(_1756_),
    .D(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__nand2_1 _5332_ (.A(_0405_),
    .B(_0889_),
    .Y(_1761_));
 sky130_fd_sc_hd__nand2_1 _5333_ (.A(_0409_),
    .B(_0456_),
    .Y(_1762_));
 sky130_fd_sc_hd__or2_1 _5334_ (.A(_3153_),
    .B(_0414_),
    .X(_1763_));
 sky130_fd_sc_hd__o2111a_1 _5335_ (.A1(_1017_),
    .A2(_0402_),
    .B1(_1761_),
    .C1(_1762_),
    .D1(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__nand2_1 _5336_ (.A(_0422_),
    .B(_3161_),
    .Y(_1765_));
 sky130_fd_sc_hd__nand2_1 _5337_ (.A(_0426_),
    .B(_3148_),
    .Y(_1766_));
 sky130_fd_sc_hd__or2_1 _5338_ (.A(_0790_),
    .B(_0431_),
    .X(_1767_));
 sky130_fd_sc_hd__o2111a_1 _5339_ (.A1(_1070_),
    .A2(_0419_),
    .B1(_1765_),
    .C1(_1766_),
    .D1(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__nand2_1 _5340_ (.A(_0447_),
    .B(_0427_),
    .Y(_1769_));
 sky130_fd_sc_hd__o21ai_1 _5341_ (.A1(_0429_),
    .A2(_0444_),
    .B1(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__a221oi_1 _5342_ (.A1(_0729_),
    .A2(_0437_),
    .B1(_0452_),
    .B2(_0441_),
    .C1(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__nand2_1 _5343_ (.A(_0465_),
    .B(_0632_),
    .Y(_1772_));
 sky130_fd_sc_hd__o21ai_1 _5344_ (.A1(_3123_),
    .A2(_0462_),
    .B1(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__a221oi_1 _5345_ (.A1(_0630_),
    .A2(_0455_),
    .B1(_3181_),
    .B2(_0459_),
    .C1(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__and4_1 _5346_ (.A(_1764_),
    .B(_1768_),
    .C(_1771_),
    .D(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__and2_1 _5347_ (.A(_1760_),
    .B(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__inv_2 _5348_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_1777_));
 sky130_fd_sc_hd__nand2_1 _5349_ (.A(_0479_),
    .B(_0707_),
    .Y(_1778_));
 sky130_fd_sc_hd__a22o_1 _5350_ (.A1(_0483_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .B1(_0485_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_1779_));
 sky130_fd_sc_hd__inv_2 _5351_ (.A(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__o211a_1 _5352_ (.A1(_1777_),
    .A2(_0476_),
    .B1(_1778_),
    .C1(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__nand2_1 _5353_ (.A(_0503_),
    .B(_0544_),
    .Y(_1782_));
 sky130_fd_sc_hd__o21ai_1 _5354_ (.A1(_1031_),
    .A2(_0500_),
    .B1(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__a221oi_1 _5355_ (.A1(_0480_),
    .A2(_0492_),
    .B1(_0745_),
    .B2(_0496_),
    .C1(_1783_),
    .Y(_1784_));
 sky130_fd_sc_hd__nand2_1 _5356_ (.A(_0514_),
    .B(_0532_),
    .Y(_1785_));
 sky130_fd_sc_hd__nand2_1 _5357_ (.A(_0519_),
    .B(_0539_),
    .Y(_1786_));
 sky130_fd_sc_hd__or2_1 _5358_ (.A(_1409_),
    .B(_0525_),
    .X(_1787_));
 sky130_fd_sc_hd__o2111a_1 _5359_ (.A1(_1655_),
    .A2(_0511_),
    .B1(_1785_),
    .C1(_1786_),
    .D1(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__nand2_1 _5360_ (.A(_0538_),
    .B(_0357_),
    .Y(_1789_));
 sky130_fd_sc_hd__nand2_1 _5361_ (.A(_0543_),
    .B(_0865_),
    .Y(_1790_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(_1789_),
    .B(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__a221oi_1 _5363_ (.A1(_0360_),
    .A2(_0531_),
    .B1(_0344_),
    .B2(_0535_),
    .C1(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__and4_1 _5364_ (.A(_1781_),
    .B(_1784_),
    .C(_1788_),
    .D(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__nand2_1 _5365_ (.A(_0557_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1794_));
 sky130_fd_sc_hd__nand2_1 _5366_ (.A(_0562_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1795_));
 sky130_fd_sc_hd__or2_1 _5367_ (.A(_1058_),
    .B(_0567_),
    .X(_1796_));
 sky130_fd_sc_hd__o2111a_1 _5368_ (.A1(_0778_),
    .A2(_0554_),
    .B1(_1794_),
    .C1(_1795_),
    .D1(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__nand2_1 _5369_ (.A(_0575_),
    .B(_0504_),
    .Y(_1798_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_0579_),
    .B(_0493_),
    .Y(_1799_));
 sky130_fd_sc_hd__or2_1 _5371_ (.A(_0498_),
    .B(_0583_),
    .X(_1800_));
 sky130_fd_sc_hd__o2111a_1 _5372_ (.A1(_0901_),
    .A2(_0572_),
    .B1(_1798_),
    .C1(_1799_),
    .D1(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__or2_1 _5373_ (.A(_0605_),
    .B(_0596_),
    .X(_1802_));
 sky130_fd_sc_hd__o221a_1 _5374_ (.A1(_0570_),
    .A2(_0589_),
    .B1(_0772_),
    .B2(_0592_),
    .C1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__o22ai_1 _5375_ (.A1(_0523_),
    .A2(_0607_),
    .B1(_0756_),
    .B2(_0610_),
    .Y(_1804_));
 sky130_fd_sc_hd__a221oi_1 _5376_ (.A1(_0508_),
    .A2(_0601_),
    .B1(_0471_),
    .B2(_0604_),
    .C1(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__and4_1 _5377_ (.A(_1797_),
    .B(_1801_),
    .C(_1803_),
    .D(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__and3_1 _5378_ (.A(_1776_),
    .B(_1793_),
    .C(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__nand2_1 _5379_ (.A(_0618_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1808_));
 sky130_fd_sc_hd__nand3_1 _5380_ (.A(_1745_),
    .B(_1807_),
    .C(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__inv_2 _5381_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_1810_));
 sky130_fd_sc_hd__a21oi_1 _5382_ (.A1(_1810_),
    .A2(_3102_),
    .B1(_2985_),
    .Y(_1811_));
 sky130_fd_sc_hd__o21a_1 _5383_ (.A1(_3103_),
    .A2(_1809_),
    .B1(_1811_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _5384_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1812_));
 sky130_fd_sc_hd__o22ai_1 _5385_ (.A1(_1690_),
    .A2(_3129_),
    .B1(_1812_),
    .B2(_3137_),
    .Y(_1813_));
 sky130_fd_sc_hd__a221oi_1 _5386_ (.A1(_0663_),
    .A2(_3114_),
    .B1(_0824_),
    .B2(_3121_),
    .C1(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__nand2_1 _5387_ (.A(_3159_),
    .B(_3116_),
    .Y(_1815_));
 sky130_fd_sc_hd__o21ai_1 _5388_ (.A1(_0623_),
    .A2(_3155_),
    .B1(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__a221oi_2 _5389_ (.A1(_3209_),
    .A2(_3146_),
    .B1(_3203_),
    .B2(_3151_),
    .C1(_1816_),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(_3173_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1818_));
 sky130_fd_sc_hd__nand2_1 _5391_ (.A(_3179_),
    .B(_0637_),
    .Y(_1819_));
 sky130_fd_sc_hd__or2_1 _5392_ (.A(_1320_),
    .B(_3186_),
    .X(_1820_));
 sky130_fd_sc_hd__o2111a_1 _5393_ (.A1(_1568_),
    .A2(_3168_),
    .B1(_1818_),
    .C1(_1819_),
    .D1(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__nand2_1 _5394_ (.A(_3201_),
    .B(_3323_),
    .Y(_1822_));
 sky130_fd_sc_hd__nand2_1 _5395_ (.A(_3207_),
    .B(_0967_),
    .Y(_1823_));
 sky130_fd_sc_hd__nand2_1 _5396_ (.A(_1822_),
    .B(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__a221oi_1 _5397_ (.A1(_0670_),
    .A2(_3193_),
    .B1(_0831_),
    .B2(_3197_),
    .C1(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__and4_1 _5398_ (.A(_1814_),
    .B(_1817_),
    .C(_1821_),
    .D(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__o22ai_1 _5399_ (.A1(_0653_),
    .A2(_3223_),
    .B1(_0815_),
    .B2(_3226_),
    .Y(_1827_));
 sky130_fd_sc_hd__a221oi_1 _5400_ (.A1(_0619_),
    .A2(_3217_),
    .B1(_0783_),
    .B2(_3220_),
    .C1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand2_1 _5401_ (.A(_3240_),
    .B(_0563_),
    .Y(_1829_));
 sky130_fd_sc_hd__o21ai_1 _5402_ (.A1(_0550_),
    .A2(_3237_),
    .B1(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__a221oi_1 _5403_ (.A1(_0586_),
    .A2(_3231_),
    .B1(_0593_),
    .B2(_3234_),
    .C1(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(_3255_),
    .B(_3087_),
    .Y(_1832_));
 sky130_fd_sc_hd__o21ai_1 _5405_ (.A1(_1210_),
    .A2(_3252_),
    .B1(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__a221oi_1 _5406_ (.A1(_3090_),
    .A2(_3246_),
    .B1(_3093_),
    .B2(_3249_),
    .C1(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__o22ai_1 _5407_ (.A1(_0764_),
    .A2(_3267_),
    .B1(_0565_),
    .B2(_3270_),
    .Y(_1835_));
 sky130_fd_sc_hd__a221oi_1 _5408_ (.A1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .A2(_3261_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .B2(_3264_),
    .C1(_1835_),
    .Y(_1836_));
 sky130_fd_sc_hd__and4_1 _5409_ (.A(_1828_),
    .B(_1831_),
    .C(_1834_),
    .D(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__o22ai_1 _5410_ (.A1(_1232_),
    .A2(_3287_),
    .B1(_1356_),
    .B2(_3290_),
    .Y(_1838_));
 sky130_fd_sc_hd__a221oi_1 _5411_ (.A1(_3391_),
    .A2(_3280_),
    .B1(_0686_),
    .B2(_3284_),
    .C1(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__nand2_1 _5412_ (.A(_3295_),
    .B(_3282_),
    .Y(_1840_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(_3299_),
    .B(_0819_),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _5414_ (.A(_3304_),
    .B(_3275_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _5415_ (.A(_3308_),
    .B(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_1843_));
 sky130_fd_sc_hd__and4_1 _5416_ (.A(_1840_),
    .B(_1841_),
    .C(_1842_),
    .D(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__o22ai_1 _5417_ (.A1(_0673_),
    .A2(_3313_),
    .B1(_0834_),
    .B2(_3316_),
    .Y(_1845_));
 sky130_fd_sc_hd__a22o_1 _5418_ (.A1(_3319_),
    .A2(_3366_),
    .B1(_3321_),
    .B2(_3370_),
    .X(_1846_));
 sky130_fd_sc_hd__nor2_1 _5419_ (.A(_1845_),
    .B(_1846_),
    .Y(_1847_));
 sky130_fd_sc_hd__o22ai_1 _5420_ (.A1(_0690_),
    .A2(_3335_),
    .B1(_3385_),
    .B2(_3338_),
    .Y(_1848_));
 sky130_fd_sc_hd__a221oi_1 _5421_ (.A1(_3362_),
    .A2(_3328_),
    .B1(_3357_),
    .B2(_3332_),
    .C1(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__and4_1 _5422_ (.A(_1839_),
    .B(_1844_),
    .C(_1847_),
    .D(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__nand2_1 _5423_ (.A(_3355_),
    .B(_3062_),
    .Y(_1851_));
 sky130_fd_sc_hd__nand2_1 _5424_ (.A(_3360_),
    .B(_3059_),
    .Y(_1852_));
 sky130_fd_sc_hd__nand2_1 _5425_ (.A(_1851_),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__a221oi_1 _5426_ (.A1(_3065_),
    .A2(_3348_),
    .B1(_3068_),
    .B2(_3352_),
    .C1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_3374_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1855_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_3379_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1856_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1855_),
    .B(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__a221oi_1 _5430_ (.A1(_3343_),
    .A2(_3368_),
    .B1(_3350_),
    .B2(_3371_),
    .C1(_1857_),
    .Y(_1858_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1859_));
 sky130_fd_sc_hd__nand2_1 _5432_ (.A(_3394_),
    .B(_3044_),
    .Y(_1860_));
 sky130_fd_sc_hd__or2_1 _5433_ (.A(_3411_),
    .B(_3399_),
    .X(_1861_));
 sky130_fd_sc_hd__o2111a_1 _5434_ (.A1(_0649_),
    .A2(_3386_),
    .B1(_1859_),
    .C1(_1860_),
    .D1(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__nand2_1 _5435_ (.A(_3415_),
    .B(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1863_));
 sky130_fd_sc_hd__o21ai_1 _5436_ (.A1(_1083_),
    .A2(_3412_),
    .B1(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__a221oi_1 _5437_ (.A1(_3071_),
    .A2(_3405_),
    .B1(_3074_),
    .B2(_3409_),
    .C1(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__and4_1 _5438_ (.A(_1854_),
    .B(_1858_),
    .C(_1862_),
    .D(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__and4_1 _5439_ (.A(_1826_),
    .B(_1837_),
    .C(_1850_),
    .D(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(_0337_),
    .B(_0438_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(_0342_),
    .B(_0434_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__a221oi_1 _5443_ (.A1(_0410_),
    .A2(_0330_),
    .B1(_0722_),
    .B2(_0334_),
    .C1(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__o22ai_1 _5444_ (.A1(_1750_),
    .A2(_0349_),
    .B1(_0389_),
    .B2(_0352_),
    .Y(_1872_));
 sky130_fd_sc_hd__a22o_1 _5445_ (.A1(_0355_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .B1(_0358_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_1873_));
 sky130_fd_sc_hd__nor2_1 _5446_ (.A(_1872_),
    .B(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__nand2_1 _5447_ (.A(_0375_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1875_));
 sky130_fd_sc_hd__o21ai_1 _5448_ (.A1(_1506_),
    .A2(_0372_),
    .B1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__a221oi_1 _5449_ (.A1(_0326_),
    .A2(_0365_),
    .B1(_0332_),
    .B2(_0369_),
    .C1(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _5450_ (.A(_0393_),
    .B(_0874_),
    .Y(_1878_));
 sky130_fd_sc_hd__o21ai_1 _5451_ (.A1(_0429_),
    .A2(_0390_),
    .B1(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__a221oi_1 _5452_ (.A1(_0876_),
    .A2(_0383_),
    .B1(_0720_),
    .B2(_0387_),
    .C1(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__and4_1 _5453_ (.A(_1871_),
    .B(_1874_),
    .C(_1877_),
    .D(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__nand2_1 _5454_ (.A(_0404_),
    .B(_0890_),
    .Y(_1882_));
 sky130_fd_sc_hd__nand2_1 _5455_ (.A(_0408_),
    .B(_0738_),
    .Y(_1883_));
 sky130_fd_sc_hd__or2_1 _5456_ (.A(_0626_),
    .B(_0413_),
    .X(_1884_));
 sky130_fd_sc_hd__o2111a_1 _5457_ (.A1(_0460_),
    .A2(_0401_),
    .B1(_1882_),
    .C1(_1883_),
    .D1(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_0421_),
    .B(_3141_),
    .Y(_1886_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_0425_),
    .B(_3175_),
    .Y(_1887_));
 sky130_fd_sc_hd__or2_1 _5460_ (.A(_0937_),
    .B(_0430_),
    .X(_1888_));
 sky130_fd_sc_hd__o2111a_1 _5461_ (.A1(_3183_),
    .A2(_0418_),
    .B1(_1886_),
    .C1(_1887_),
    .D1(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__nand2_1 _5462_ (.A(_0446_),
    .B(_0729_),
    .Y(_1890_));
 sky130_fd_sc_hd__o21ai_1 _5463_ (.A1(_0731_),
    .A2(_0443_),
    .B1(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__a221oi_1 _5464_ (.A1(_0452_),
    .A2(_0436_),
    .B1(_0456_),
    .B2(_0440_),
    .C1(_1891_),
    .Y(_1892_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_0464_),
    .B(_0795_),
    .Y(_1893_));
 sky130_fd_sc_hd__o21ai_1 _5466_ (.A1(_3132_),
    .A2(_0461_),
    .B1(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__a221oi_1 _5467_ (.A1(_3181_),
    .A2(_0454_),
    .B1(_0632_),
    .B2(_0458_),
    .C1(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__and4_1 _5468_ (.A(_1885_),
    .B(_1889_),
    .C(_1892_),
    .D(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__and2_1 _5469_ (.A(_1881_),
    .B(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__nand2_1 _5470_ (.A(_0478_),
    .B(_0377_),
    .Y(_1898_));
 sky130_fd_sc_hd__a22o_1 _5471_ (.A1(_0482_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .B1(_0484_),
    .B2(_0865_),
    .X(_1899_));
 sky130_fd_sc_hd__inv_2 _5472_ (.A(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__o211a_1 _5473_ (.A1(_0371_),
    .A2(_0475_),
    .B1(_1898_),
    .C1(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__nand2_1 _5474_ (.A(_0502_),
    .B(_0539_),
    .Y(_1902_));
 sky130_fd_sc_hd__o21ai_1 _5475_ (.A1(_1159_),
    .A2(_0499_),
    .B1(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__a221oi_1 _5476_ (.A1(_0745_),
    .A2(_0491_),
    .B1(_0486_),
    .B2(_0495_),
    .C1(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__nand2_1 _5477_ (.A(_0513_),
    .B(_0363_),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _5478_ (.A(_0518_),
    .B(_0528_),
    .Y(_1906_));
 sky130_fd_sc_hd__or2_1 _5479_ (.A(_1533_),
    .B(_0524_),
    .X(_1907_));
 sky130_fd_sc_hd__o2111a_1 _5480_ (.A1(_1777_),
    .A2(_0510_),
    .B1(_1905_),
    .C1(_1906_),
    .D1(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__nand2_1 _5481_ (.A(_0537_),
    .B(_0360_),
    .Y(_1909_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_0542_),
    .B(_0357_),
    .Y(_1910_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_1909_),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__a221oi_1 _5484_ (.A1(_0344_),
    .A2(_0530_),
    .B1(_0339_),
    .B2(_0534_),
    .C1(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__and4_1 _5485_ (.A(_1901_),
    .B(_1904_),
    .C(_1908_),
    .D(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__nand2_1 _5486_ (.A(_0556_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1915_));
 sky130_fd_sc_hd__or2_1 _5488_ (.A(_1186_),
    .B(_0566_),
    .X(_1916_));
 sky130_fd_sc_hd__o2111a_1 _5489_ (.A1(_0924_),
    .A2(_0553_),
    .B1(_1914_),
    .C1(_1915_),
    .D1(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__nand2_1 _5490_ (.A(_0574_),
    .B(_0520_),
    .Y(_1918_));
 sky130_fd_sc_hd__nand2_1 _5491_ (.A(_0578_),
    .B(_0497_),
    .Y(_1919_));
 sky130_fd_sc_hd__or2_1 _5492_ (.A(_0750_),
    .B(_0582_),
    .X(_1920_));
 sky130_fd_sc_hd__o2111a_1 _5493_ (.A1(_0523_),
    .A2(_0571_),
    .B1(_1918_),
    .C1(_1919_),
    .D1(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__or2_1 _5494_ (.A(_0608_),
    .B(_0595_),
    .X(_1922_));
 sky130_fd_sc_hd__o221a_1 _5495_ (.A1(_0605_),
    .A2(_0588_),
    .B1(_0570_),
    .B2(_0591_),
    .C1(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__o22ai_1 _5496_ (.A1(_0756_),
    .A2(_0606_),
    .B1(_0509_),
    .B2(_0609_),
    .Y(_1924_));
 sky130_fd_sc_hd__a221oi_2 _5497_ (.A1(_0471_),
    .A2(_0600_),
    .B1(_0480_),
    .B2(_0603_),
    .C1(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__and4_1 _5498_ (.A(_1917_),
    .B(_1921_),
    .C(_1923_),
    .D(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__and3_1 _5499_ (.A(_1897_),
    .B(_1913_),
    .C(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__nand2_1 _5500_ (.A(_0617_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1928_));
 sky130_fd_sc_hd__nand3_1 _5501_ (.A(_1867_),
    .B(_1927_),
    .C(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__inv_2 _5502_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_1930_));
 sky130_fd_sc_hd__a21oi_1 _5503_ (.A1(_1930_),
    .A2(_3102_),
    .B1(_2984_),
    .Y(_1931_));
 sky130_fd_sc_hd__o21a_1 _5504_ (.A1(_0932_),
    .A2(_1929_),
    .B1(_1931_),
    .X(_0287_));
 sky130_fd_sc_hd__o22ai_1 _5505_ (.A1(_1812_),
    .A2(_3129_),
    .B1(_3312_),
    .B2(_3137_),
    .Y(_1932_));
 sky130_fd_sc_hd__a221oi_1 _5506_ (.A1(_0824_),
    .A2(_3114_),
    .B1(_0967_),
    .B2(_3121_),
    .C1(_1932_),
    .Y(_1933_));
 sky130_fd_sc_hd__nand2_1 _5507_ (.A(_3159_),
    .B(_3209_),
    .Y(_1934_));
 sky130_fd_sc_hd__o21ai_1 _5508_ (.A1(_0787_),
    .A2(_3155_),
    .B1(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__a221oi_1 _5509_ (.A1(_3203_),
    .A2(_3146_),
    .B1(_3190_),
    .B2(_3151_),
    .C1(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _5510_ (.A(_3173_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _5511_ (.A(_3179_),
    .B(_0799_),
    .Y(_1938_));
 sky130_fd_sc_hd__or2_1 _5512_ (.A(_1444_),
    .B(_3186_),
    .X(_1939_));
 sky130_fd_sc_hd__o2111a_1 _5513_ (.A1(_1690_),
    .A2(_3168_),
    .B1(_1937_),
    .C1(_1938_),
    .D1(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__nand2_1 _5514_ (.A(_3201_),
    .B(_0670_),
    .Y(_1941_));
 sky130_fd_sc_hd__nand2_1 _5515_ (.A(_3207_),
    .B(_3323_),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5516_ (.A(_1941_),
    .B(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__a221oi_1 _5517_ (.A1(_0831_),
    .A2(_3193_),
    .B1(_3275_),
    .B2(_3197_),
    .C1(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__and4_1 _5518_ (.A(_1933_),
    .B(_1936_),
    .C(_1940_),
    .D(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__o22ai_1 _5519_ (.A1(_0815_),
    .A2(_3223_),
    .B1(_0960_),
    .B2(_3226_),
    .Y(_1946_));
 sky130_fd_sc_hd__a221oi_1 _5520_ (.A1(_0783_),
    .A2(_3217_),
    .B1(_0586_),
    .B2(_3220_),
    .C1(_1946_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _5521_ (.A(_3240_),
    .B(_0549_),
    .Y(_1948_));
 sky130_fd_sc_hd__o21ai_1 _5522_ (.A1(_0764_),
    .A2(_3237_),
    .B1(_1948_),
    .Y(_1949_));
 sky130_fd_sc_hd__a221oi_1 _5523_ (.A1(_0593_),
    .A2(_3231_),
    .B1(_0563_),
    .B2(_3234_),
    .C1(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _5524_ (.A(_3255_),
    .B(_3090_),
    .Y(_1951_));
 sky130_fd_sc_hd__o21ai_1 _5525_ (.A1(_3236_),
    .A2(_3252_),
    .B1(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__a221oi_1 _5526_ (.A1(_3093_),
    .A2(_3246_),
    .B1(_3096_),
    .B2(_3249_),
    .C1(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__o22ai_1 _5527_ (.A1(_0565_),
    .A2(_3267_),
    .B1(_0767_),
    .B2(_3270_),
    .Y(_1954_));
 sky130_fd_sc_hd__a221oi_1 _5528_ (.A1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .A2(_3261_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .B2(_3264_),
    .C1(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__and4_1 _5529_ (.A(_1947_),
    .B(_1950_),
    .C(_1953_),
    .D(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__o22ai_1 _5530_ (.A1(_1356_),
    .A2(_3287_),
    .B1(_1480_),
    .B2(_3290_),
    .Y(_1957_));
 sky130_fd_sc_hd__a221oi_1 _5531_ (.A1(_0686_),
    .A2(_3280_),
    .B1(_3396_),
    .B2(_3284_),
    .C1(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__nand2_1 _5532_ (.A(_3295_),
    .B(_0657_),
    .Y(_1959_));
 sky130_fd_sc_hd__nand2_1 _5533_ (.A(_3299_),
    .B(_3326_),
    .Y(_1960_));
 sky130_fd_sc_hd__nand2_1 _5534_ (.A(_3304_),
    .B(_3282_),
    .Y(_1961_));
 sky130_fd_sc_hd__nand2_1 _5535_ (.A(_3308_),
    .B(_0819_),
    .Y(_1962_));
 sky130_fd_sc_hd__and4_1 _5536_ (.A(_1959_),
    .B(_1960_),
    .C(_1961_),
    .D(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__o22ai_1 _5537_ (.A1(_0834_),
    .A2(_3313_),
    .B1(_0975_),
    .B2(_3316_),
    .Y(_1964_));
 sky130_fd_sc_hd__a22o_1 _5538_ (.A1(_3319_),
    .A2(_3370_),
    .B1(_3321_),
    .B2(_3381_),
    .X(_1965_));
 sky130_fd_sc_hd__nor2_1 _5539_ (.A(_1964_),
    .B(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__o22ai_1 _5540_ (.A1(_3385_),
    .A2(_3335_),
    .B1(_0685_),
    .B2(_3338_),
    .Y(_1967_));
 sky130_fd_sc_hd__a221oi_1 _5541_ (.A1(_3357_),
    .A2(_3328_),
    .B1(_3343_),
    .B2(_3332_),
    .C1(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__and4_1 _5542_ (.A(_1958_),
    .B(_1963_),
    .C(_1966_),
    .D(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__nand2_1 _5543_ (.A(_3355_),
    .B(_3065_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _5544_ (.A(_3360_),
    .B(_3062_),
    .Y(_1971_));
 sky130_fd_sc_hd__nand2_1 _5545_ (.A(_1970_),
    .B(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__a221oi_1 _5546_ (.A1(_3068_),
    .A2(_3348_),
    .B1(_3071_),
    .B2(_3352_),
    .C1(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__nand2_1 _5547_ (.A(_3374_),
    .B(_0693_),
    .Y(_1974_));
 sky130_fd_sc_hd__nand2_1 _5548_ (.A(_3379_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2_1 _5549_ (.A(_1974_),
    .B(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__a221oi_1 _5550_ (.A1(_3350_),
    .A2(_3368_),
    .B1(_3403_),
    .B2(_3371_),
    .C1(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _5551_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_1978_));
 sky130_fd_sc_hd__nand2_1 _5552_ (.A(_3394_),
    .B(_3056_),
    .Y(_1979_));
 sky130_fd_sc_hd__or2_1 _5553_ (.A(_3251_),
    .B(_3399_),
    .X(_1980_));
 sky130_fd_sc_hd__o2111a_1 _5554_ (.A1(_0811_),
    .A2(_3386_),
    .B1(_1978_),
    .C1(_1979_),
    .D1(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__nand2_1 _5555_ (.A(_3415_),
    .B(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1982_));
 sky130_fd_sc_hd__o21ai_1 _5556_ (.A1(_1210_),
    .A2(_3412_),
    .B1(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__a221oi_1 _5557_ (.A1(_3074_),
    .A2(_3405_),
    .B1(_3078_),
    .B2(_3409_),
    .C1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__and4_1 _5558_ (.A(_1973_),
    .B(_1977_),
    .C(_1981_),
    .D(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__and4_1 _5559_ (.A(_1945_),
    .B(_1956_),
    .C(_1969_),
    .D(_1985_),
    .X(_1986_));
 sky130_fd_sc_hd__nand2_1 _5560_ (.A(_0337_),
    .B(_0410_),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _5561_ (.A(_0342_),
    .B(_0438_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5562_ (.A(_1987_),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__a221oi_1 _5563_ (.A1(_0722_),
    .A2(_0330_),
    .B1(_0876_),
    .B2(_0334_),
    .C1(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__o22ai_1 _5564_ (.A1(_0389_),
    .A2(_0349_),
    .B1(_0442_),
    .B2(_0352_),
    .Y(_1991_));
 sky130_fd_sc_hd__a22o_1 _5565_ (.A1(_0355_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .B1(_0358_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_1992_));
 sky130_fd_sc_hd__nor2_1 _5566_ (.A(_1991_),
    .B(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__nand2_1 _5567_ (.A(_0375_),
    .B(_0713_),
    .Y(_1994_));
 sky130_fd_sc_hd__o21ai_1 _5568_ (.A1(_1628_),
    .A2(_0372_),
    .B1(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__a221oi_1 _5569_ (.A1(_0332_),
    .A2(_0365_),
    .B1(_0381_),
    .B2(_0369_),
    .C1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_1 _5570_ (.A(_0393_),
    .B(_1012_),
    .Y(_1997_));
 sky130_fd_sc_hd__o21ai_1 _5571_ (.A1(_0731_),
    .A2(_0390_),
    .B1(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__a221oi_1 _5572_ (.A1(_0720_),
    .A2(_0383_),
    .B1(_0874_),
    .B2(_0387_),
    .C1(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__and4_1 _5573_ (.A(_1990_),
    .B(_1993_),
    .C(_1996_),
    .D(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(_0404_),
    .B(_3161_),
    .Y(_2001_));
 sky130_fd_sc_hd__nand2_1 _5575_ (.A(_0408_),
    .B(_0889_),
    .Y(_2002_));
 sky130_fd_sc_hd__or2_1 _5576_ (.A(_0790_),
    .B(_0413_),
    .X(_2003_));
 sky130_fd_sc_hd__o2111a_1 _5577_ (.A1(_3153_),
    .A2(_0401_),
    .B1(_2001_),
    .C1(_2002_),
    .D1(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__nand2_1 _5578_ (.A(_0421_),
    .B(_3148_),
    .Y(_2005_));
 sky130_fd_sc_hd__nand2_1 _5579_ (.A(_0425_),
    .B(_0630_),
    .Y(_2006_));
 sky130_fd_sc_hd__or2_1 _5580_ (.A(_1070_),
    .B(_0430_),
    .X(_2007_));
 sky130_fd_sc_hd__o2111a_1 _5581_ (.A1(_0634_),
    .A2(_0418_),
    .B1(_2005_),
    .C1(_2006_),
    .D1(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__nand2_1 _5582_ (.A(_0446_),
    .B(_0452_),
    .Y(_2009_));
 sky130_fd_sc_hd__o21ai_1 _5583_ (.A1(_0417_),
    .A2(_0443_),
    .B1(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__a221oi_1 _5584_ (.A1(_0456_),
    .A2(_0436_),
    .B1(_0738_),
    .B2(_0440_),
    .C1(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _5585_ (.A(_0464_),
    .B(_3131_),
    .Y(_2012_));
 sky130_fd_sc_hd__o21ai_1 _5586_ (.A1(_0623_),
    .A2(_0461_),
    .B1(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hd__a221oi_1 _5587_ (.A1(_0632_),
    .A2(_0454_),
    .B1(_0795_),
    .B2(_0458_),
    .C1(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__and4_1 _5588_ (.A(_2004_),
    .B(_2008_),
    .C(_2011_),
    .D(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__and2_1 _5589_ (.A(_2000_),
    .B(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__nand2_1 _5590_ (.A(_0478_),
    .B(_0709_),
    .Y(_2017_));
 sky130_fd_sc_hd__a22o_1 _5591_ (.A1(_0482_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .B1(_0484_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_2018_));
 sky130_fd_sc_hd__inv_2 _5592_ (.A(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__o211a_1 _5593_ (.A1(_0708_),
    .A2(_0475_),
    .B1(_2017_),
    .C1(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__nand2_1 _5594_ (.A(_0502_),
    .B(_0528_),
    .Y(_2021_));
 sky130_fd_sc_hd__o21ai_1 _5595_ (.A1(_1285_),
    .A2(_0499_),
    .B1(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__a221oi_1 _5596_ (.A1(_0486_),
    .A2(_0491_),
    .B1(_0544_),
    .B2(_0495_),
    .C1(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2_1 _5597_ (.A(_0513_),
    .B(_0367_),
    .Y(_2024_));
 sky130_fd_sc_hd__nand2_1 _5598_ (.A(_0518_),
    .B(_0532_),
    .Y(_2025_));
 sky130_fd_sc_hd__or2_1 _5599_ (.A(_1655_),
    .B(_0524_),
    .X(_2026_));
 sky130_fd_sc_hd__o2111a_1 _5600_ (.A1(_0371_),
    .A2(_0510_),
    .B1(_2024_),
    .C1(_2025_),
    .D1(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(_0537_),
    .B(_0344_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_0542_),
    .B(_0360_),
    .Y(_2029_));
 sky130_fd_sc_hd__nand2_1 _5603_ (.A(_2028_),
    .B(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__a221oi_1 _5604_ (.A1(_0339_),
    .A2(_0530_),
    .B1(_0326_),
    .B2(_0534_),
    .C1(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__and4_1 _5605_ (.A(_2020_),
    .B(_2023_),
    .C(_2027_),
    .D(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_0556_),
    .B(_0493_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand2_1 _5607_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_2034_));
 sky130_fd_sc_hd__or2_1 _5608_ (.A(_0498_),
    .B(_0566_),
    .X(_2035_));
 sky130_fd_sc_hd__o2111a_1 _5609_ (.A1(_1058_),
    .A2(_0553_),
    .B1(_2033_),
    .C1(_2034_),
    .D1(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(_0574_),
    .B(_0522_),
    .Y(_2037_));
 sky130_fd_sc_hd__nand2_1 _5611_ (.A(_0578_),
    .B(_0504_),
    .Y(_2038_));
 sky130_fd_sc_hd__or2_1 _5612_ (.A(_0901_),
    .B(_0582_),
    .X(_2039_));
 sky130_fd_sc_hd__o2111a_1 _5613_ (.A1(_0756_),
    .A2(_0571_),
    .B1(_2037_),
    .C1(_2038_),
    .D1(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__or2_1 _5614_ (.A(_0778_),
    .B(_0595_),
    .X(_2041_));
 sky130_fd_sc_hd__o221a_1 _5615_ (.A1(_0608_),
    .A2(_0588_),
    .B1(_0605_),
    .B2(_0591_),
    .C1(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__o22ai_1 _5616_ (.A1(_0509_),
    .A2(_0606_),
    .B1(_0472_),
    .B2(_0609_),
    .Y(_2043_));
 sky130_fd_sc_hd__a221oi_1 _5617_ (.A1(_0480_),
    .A2(_0600_),
    .B1(_0745_),
    .B2(_0603_),
    .C1(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__and4_1 _5618_ (.A(_2036_),
    .B(_2040_),
    .C(_2042_),
    .D(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__and3_1 _5619_ (.A(_2016_),
    .B(_2032_),
    .C(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__nand2_1 _5620_ (.A(_0617_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_2047_));
 sky130_fd_sc_hd__nand3_1 _5621_ (.A(_1986_),
    .B(_2046_),
    .C(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__inv_2 _5622_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2049_));
 sky130_fd_sc_hd__a21oi_1 _5623_ (.A1(_2049_),
    .A2(_3102_),
    .B1(_2984_),
    .Y(_2050_));
 sky130_fd_sc_hd__o21a_1 _5624_ (.A1(_0932_),
    .A2(_2048_),
    .B1(_2050_),
    .X(_0286_));
 sky130_fd_sc_hd__o22ai_1 _5625_ (.A1(_3312_),
    .A2(_3129_),
    .B1(_3315_),
    .B2(_3137_),
    .Y(_2051_));
 sky130_fd_sc_hd__a221oi_1 _5626_ (.A1(_0967_),
    .A2(_3114_),
    .B1(_3323_),
    .B2(_3121_),
    .C1(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__nand2_1 _5627_ (.A(_3159_),
    .B(_3203_),
    .Y(_2053_));
 sky130_fd_sc_hd__o21ai_1 _5628_ (.A1(_0934_),
    .A2(_3155_),
    .B1(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__a221oi_1 _5629_ (.A1(_3190_),
    .A2(_3146_),
    .B1(_3195_),
    .B2(_3151_),
    .C1(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__nand2_1 _5630_ (.A(_3173_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _5631_ (.A(_3179_),
    .B(_0661_),
    .Y(_2057_));
 sky130_fd_sc_hd__or2_1 _5632_ (.A(_1568_),
    .B(_3186_),
    .X(_2058_));
 sky130_fd_sc_hd__o2111a_1 _5633_ (.A1(_1812_),
    .A2(_3168_),
    .B1(_2056_),
    .C1(_2057_),
    .D1(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(_3201_),
    .B(_0831_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _5635_ (.A(_3207_),
    .B(_0670_),
    .Y(_2061_));
 sky130_fd_sc_hd__nand2_1 _5636_ (.A(_2060_),
    .B(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__a221oi_1 _5637_ (.A1(_3275_),
    .A2(_3193_),
    .B1(_3282_),
    .B2(_3197_),
    .C1(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__and4_1 _5638_ (.A(_2052_),
    .B(_2055_),
    .C(_2059_),
    .D(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__o22ai_1 _5639_ (.A1(_0960_),
    .A2(_3223_),
    .B1(_0590_),
    .B2(_3226_),
    .Y(_2065_));
 sky130_fd_sc_hd__a221oi_1 _5640_ (.A1(_0586_),
    .A2(_3217_),
    .B1(_0593_),
    .B2(_3220_),
    .C1(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__nand2_1 _5641_ (.A(_3240_),
    .B(_0558_),
    .Y(_2067_));
 sky130_fd_sc_hd__o21ai_1 _5642_ (.A1(_0565_),
    .A2(_3237_),
    .B1(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__a221oi_1 _5643_ (.A1(_0563_),
    .A2(_3231_),
    .B1(_0549_),
    .B2(_3234_),
    .C1(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__nand2_1 _5644_ (.A(_3255_),
    .B(_3093_),
    .Y(_2070_));
 sky130_fd_sc_hd__o21ai_1 _5645_ (.A1(_3266_),
    .A2(_3252_),
    .B1(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__a221oi_1 _5646_ (.A1(_3096_),
    .A2(_3246_),
    .B1(_3099_),
    .B2(_3249_),
    .C1(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__o22ai_1 _5647_ (.A1(_0767_),
    .A2(_3267_),
    .B1(_0581_),
    .B2(_3270_),
    .Y(_2073_));
 sky130_fd_sc_hd__a221oi_1 _5648_ (.A1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .A2(_3261_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .B2(_3264_),
    .C1(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__and4_1 _5649_ (.A(_2066_),
    .B(_2069_),
    .C(_2072_),
    .D(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__o22ai_1 _5650_ (.A1(_1480_),
    .A2(_3287_),
    .B1(_3398_),
    .B2(_3290_),
    .Y(_2076_));
 sky130_fd_sc_hd__a221oi_1 _5651_ (.A1(_3396_),
    .A2(_3280_),
    .B1(_0688_),
    .B2(_3284_),
    .C1(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__nand2_1 _5652_ (.A(_3295_),
    .B(_0819_),
    .Y(_2078_));
 sky130_fd_sc_hd__nand2_1 _5653_ (.A(_3299_),
    .B(_3330_),
    .Y(_2079_));
 sky130_fd_sc_hd__nand2_1 _5654_ (.A(_3304_),
    .B(_0657_),
    .Y(_2080_));
 sky130_fd_sc_hd__nand2_1 _5655_ (.A(_3308_),
    .B(_3326_),
    .Y(_2081_));
 sky130_fd_sc_hd__and4_1 _5656_ (.A(_2078_),
    .B(_2079_),
    .C(_2080_),
    .D(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__o22ai_1 _5657_ (.A1(_0975_),
    .A2(_3313_),
    .B1(_1105_),
    .B2(_3316_),
    .Y(_2083_));
 sky130_fd_sc_hd__a22o_1 _5658_ (.A1(_3319_),
    .A2(_3381_),
    .B1(_3321_),
    .B2(_3376_),
    .X(_2084_));
 sky130_fd_sc_hd__nor2_1 _5659_ (.A(_2083_),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__o22ai_1 _5660_ (.A1(_0685_),
    .A2(_3335_),
    .B1(_0846_),
    .B2(_3338_),
    .Y(_2086_));
 sky130_fd_sc_hd__a221oi_1 _5661_ (.A1(_3343_),
    .A2(_3328_),
    .B1(_3350_),
    .B2(_3332_),
    .C1(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__and4_1 _5662_ (.A(_2077_),
    .B(_2082_),
    .C(_2085_),
    .D(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__nand2_1 _5663_ (.A(_3355_),
    .B(_3068_),
    .Y(_2089_));
 sky130_fd_sc_hd__nand2_1 _5664_ (.A(_3360_),
    .B(_3065_),
    .Y(_2090_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(_2089_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__a221oi_1 _5666_ (.A1(_3071_),
    .A2(_3348_),
    .B1(_3074_),
    .B2(_3352_),
    .C1(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__nand2_1 _5667_ (.A(_3374_),
    .B(_0851_),
    .Y(_2093_));
 sky130_fd_sc_hd__nand2_1 _5668_ (.A(_3379_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_2094_));
 sky130_fd_sc_hd__nand2_1 _5669_ (.A(_2093_),
    .B(_2094_),
    .Y(_2095_));
 sky130_fd_sc_hd__a221oi_1 _5670_ (.A1(_3403_),
    .A2(_3368_),
    .B1(_3407_),
    .B2(_3371_),
    .C1(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _5671_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_2097_));
 sky130_fd_sc_hd__nand2_1 _5672_ (.A(_3394_),
    .B(_3059_),
    .Y(_2098_));
 sky130_fd_sc_hd__or2_1 _5673_ (.A(_0649_),
    .B(_3399_),
    .X(_2099_));
 sky130_fd_sc_hd__o2111a_1 _5674_ (.A1(_0956_),
    .A2(_3386_),
    .B1(_2097_),
    .C1(_2098_),
    .D1(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_3415_),
    .B(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_2101_));
 sky130_fd_sc_hd__o21ai_1 _5676_ (.A1(_3236_),
    .A2(_3412_),
    .B1(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__a221oi_1 _5677_ (.A1(_3078_),
    .A2(_3405_),
    .B1(_3081_),
    .B2(_3409_),
    .C1(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__and4_1 _5678_ (.A(_2092_),
    .B(_2096_),
    .C(_2100_),
    .D(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__and4_1 _5679_ (.A(_2064_),
    .B(_2075_),
    .C(_2088_),
    .D(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__nand2_1 _5680_ (.A(_0337_),
    .B(_0722_),
    .Y(_2106_));
 sky130_fd_sc_hd__nand2_1 _5681_ (.A(_0342_),
    .B(_0410_),
    .Y(_2107_));
 sky130_fd_sc_hd__nand2_1 _5682_ (.A(_2106_),
    .B(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__a221oi_1 _5683_ (.A1(_0876_),
    .A2(_0330_),
    .B1(_0720_),
    .B2(_0334_),
    .C1(_2108_),
    .Y(_2109_));
 sky130_fd_sc_hd__o22ai_1 _5684_ (.A1(_0442_),
    .A2(_0349_),
    .B1(_0734_),
    .B2(_0352_),
    .Y(_2110_));
 sky130_fd_sc_hd__a22o_1 _5685_ (.A1(_0355_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .B1(_0358_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_2111_));
 sky130_fd_sc_hd__nor2_1 _5686_ (.A(_2110_),
    .B(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__nand2_1 _5687_ (.A(_0375_),
    .B(_0714_),
    .Y(_2113_));
 sky130_fd_sc_hd__o21ai_1 _5688_ (.A1(_1750_),
    .A2(_0372_),
    .B1(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__a221oi_1 _5689_ (.A1(_0381_),
    .A2(_0365_),
    .B1(_0385_),
    .B2(_0369_),
    .C1(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_0393_),
    .B(_0427_),
    .Y(_2116_));
 sky130_fd_sc_hd__o21ai_1 _5691_ (.A1(_0417_),
    .A2(_0390_),
    .B1(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__a221oi_1 _5692_ (.A1(_0874_),
    .A2(_0383_),
    .B1(_1012_),
    .B2(_0387_),
    .C1(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__and4_1 _5693_ (.A(_2109_),
    .B(_2112_),
    .C(_2115_),
    .D(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__nand2_1 _5694_ (.A(_0404_),
    .B(_3141_),
    .Y(_2120_));
 sky130_fd_sc_hd__nand2_1 _5695_ (.A(_0408_),
    .B(_0890_),
    .Y(_2121_));
 sky130_fd_sc_hd__or2_1 _5696_ (.A(_0937_),
    .B(_0413_),
    .X(_2122_));
 sky130_fd_sc_hd__o2111a_1 _5697_ (.A1(_0626_),
    .A2(_0401_),
    .B1(_2120_),
    .C1(_2121_),
    .D1(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__nand2_1 _5698_ (.A(_0421_),
    .B(_3175_),
    .Y(_2124_));
 sky130_fd_sc_hd__nand2_1 _5699_ (.A(_0425_),
    .B(_3181_),
    .Y(_2125_));
 sky130_fd_sc_hd__or2_1 _5700_ (.A(_3183_),
    .B(_0430_),
    .X(_2126_));
 sky130_fd_sc_hd__o2111a_1 _5701_ (.A1(_3165_),
    .A2(_0418_),
    .B1(_2124_),
    .C1(_2125_),
    .D1(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__nand2_1 _5702_ (.A(_0446_),
    .B(_0456_),
    .Y(_2128_));
 sky130_fd_sc_hd__o21ai_1 _5703_ (.A1(_0727_),
    .A2(_0443_),
    .B1(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__a221oi_1 _5704_ (.A1(_0738_),
    .A2(_0436_),
    .B1(_0889_),
    .B2(_0440_),
    .C1(_2129_),
    .Y(_2130_));
 sky130_fd_sc_hd__nand2_1 _5705_ (.A(_0464_),
    .B(_3104_),
    .Y(_2131_));
 sky130_fd_sc_hd__o21ai_1 _5706_ (.A1(_0787_),
    .A2(_0461_),
    .B1(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__a221oi_1 _5707_ (.A1(_0795_),
    .A2(_0454_),
    .B1(_3131_),
    .B2(_0458_),
    .C1(_2132_),
    .Y(_2133_));
 sky130_fd_sc_hd__and4_1 _5708_ (.A(_2123_),
    .B(_2127_),
    .C(_2130_),
    .D(_2133_),
    .X(_2134_));
 sky130_fd_sc_hd__and2_1 _5709_ (.A(_2119_),
    .B(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__nand2_1 _5710_ (.A(_0478_),
    .B(_0865_),
    .Y(_2136_));
 sky130_fd_sc_hd__a22o_1 _5711_ (.A1(_0482_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .B1(_0484_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_2137_));
 sky130_fd_sc_hd__inv_2 _5712_ (.A(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__o211a_1 _5713_ (.A1(_0348_),
    .A2(_0475_),
    .B1(_2136_),
    .C1(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__nand2_1 _5714_ (.A(_0502_),
    .B(_0532_),
    .Y(_2140_));
 sky130_fd_sc_hd__o21ai_1 _5715_ (.A1(_1409_),
    .A2(_0499_),
    .B1(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__a221oi_1 _5716_ (.A1(_0544_),
    .A2(_0491_),
    .B1(_0539_),
    .B2(_0495_),
    .C1(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__nand2_1 _5717_ (.A(_0513_),
    .B(_0707_),
    .Y(_2143_));
 sky130_fd_sc_hd__nand2_1 _5718_ (.A(_0518_),
    .B(_0363_),
    .Y(_2144_));
 sky130_fd_sc_hd__or2_1 _5719_ (.A(_1777_),
    .B(_0524_),
    .X(_2145_));
 sky130_fd_sc_hd__o2111a_1 _5720_ (.A1(_0708_),
    .A2(_0510_),
    .B1(_2143_),
    .C1(_2144_),
    .D1(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__nand2_1 _5721_ (.A(_0537_),
    .B(_0339_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand2_1 _5722_ (.A(_0542_),
    .B(_0344_),
    .Y(_2148_));
 sky130_fd_sc_hd__nand2_1 _5723_ (.A(_2147_),
    .B(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__a221oi_1 _5724_ (.A1(_0326_),
    .A2(_0530_),
    .B1(_0332_),
    .B2(_0534_),
    .C1(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__and4_1 _5725_ (.A(_2139_),
    .B(_2142_),
    .C(_2146_),
    .D(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__nand2_1 _5726_ (.A(_0556_),
    .B(_0497_),
    .Y(_2152_));
 sky130_fd_sc_hd__nand2_1 _5727_ (.A(_0561_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_2153_));
 sky130_fd_sc_hd__or2_1 _5728_ (.A(_0750_),
    .B(_0566_),
    .X(_2154_));
 sky130_fd_sc_hd__o2111a_1 _5729_ (.A1(_1186_),
    .A2(_0553_),
    .B1(_2152_),
    .C1(_2153_),
    .D1(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__nand2_1 _5730_ (.A(_0574_),
    .B(_0515_),
    .Y(_2156_));
 sky130_fd_sc_hd__nand2_1 _5731_ (.A(_0578_),
    .B(_0520_),
    .Y(_2157_));
 sky130_fd_sc_hd__or2_1 _5732_ (.A(_0523_),
    .B(_0582_),
    .X(_2158_));
 sky130_fd_sc_hd__o2111a_1 _5733_ (.A1(_0509_),
    .A2(_0571_),
    .B1(_2156_),
    .C1(_2157_),
    .D1(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__or2_1 _5734_ (.A(_0924_),
    .B(_0595_),
    .X(_2160_));
 sky130_fd_sc_hd__o221a_1 _5735_ (.A1(_0778_),
    .A2(_0588_),
    .B1(_0608_),
    .B2(_0591_),
    .C1(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__o22ai_1 _5736_ (.A1(_0472_),
    .A2(_0606_),
    .B1(_0744_),
    .B2(_0609_),
    .Y(_2162_));
 sky130_fd_sc_hd__a221oi_1 _5737_ (.A1(_0745_),
    .A2(_0600_),
    .B1(_0486_),
    .B2(_0603_),
    .C1(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__and4_1 _5738_ (.A(_2155_),
    .B(_2159_),
    .C(_2161_),
    .D(_2163_),
    .X(_2164_));
 sky130_fd_sc_hd__and3_1 _5739_ (.A(_2135_),
    .B(_2151_),
    .C(_2164_),
    .X(_2165_));
 sky130_fd_sc_hd__nand2_1 _5740_ (.A(_0617_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_2166_));
 sky130_fd_sc_hd__nand3_1 _5741_ (.A(_2105_),
    .B(_2165_),
    .C(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__inv_2 _5742_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2168_));
 sky130_fd_sc_hd__a21oi_1 _5743_ (.A1(_2168_),
    .A2(_3102_),
    .B1(_2984_),
    .Y(_2169_));
 sky130_fd_sc_hd__o21a_1 _5744_ (.A1(_0932_),
    .A2(_2167_),
    .B1(_2169_),
    .X(_0285_));
 sky130_fd_sc_hd__o22ai_1 _5745_ (.A1(_3315_),
    .A2(_3129_),
    .B1(_0668_),
    .B2(_3137_),
    .Y(_2170_));
 sky130_fd_sc_hd__a221oi_1 _5746_ (.A1(_3323_),
    .A2(_3114_),
    .B1(_0670_),
    .B2(_3121_),
    .C1(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__nand2_1 _5747_ (.A(_3159_),
    .B(_3190_),
    .Y(_2172_));
 sky130_fd_sc_hd__o21ai_1 _5748_ (.A1(_1067_),
    .A2(_3155_),
    .B1(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__a221oi_1 _5749_ (.A1(_3195_),
    .A2(_3146_),
    .B1(_0637_),
    .B2(_3151_),
    .C1(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _5750_ (.A(_3173_),
    .B(_0799_),
    .Y(_2175_));
 sky130_fd_sc_hd__nand2_1 _5751_ (.A(_3179_),
    .B(_3301_),
    .Y(_2176_));
 sky130_fd_sc_hd__or2_1 _5752_ (.A(_1690_),
    .B(_3186_),
    .X(_2177_));
 sky130_fd_sc_hd__o2111a_1 _5753_ (.A1(_3312_),
    .A2(_3168_),
    .B1(_2175_),
    .C1(_2176_),
    .D1(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__nand2_1 _5754_ (.A(_3201_),
    .B(_3275_),
    .Y(_2179_));
 sky130_fd_sc_hd__nand2_1 _5755_ (.A(_3207_),
    .B(_0831_),
    .Y(_2180_));
 sky130_fd_sc_hd__nand2_1 _5756_ (.A(_2179_),
    .B(_2180_),
    .Y(_2181_));
 sky130_fd_sc_hd__a221oi_1 _5757_ (.A1(_3282_),
    .A2(_3193_),
    .B1(_0657_),
    .B2(_3197_),
    .C1(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__and4_1 _5758_ (.A(_2171_),
    .B(_2174_),
    .C(_2178_),
    .D(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__o22ai_1 _5759_ (.A1(_0590_),
    .A2(_3223_),
    .B1(_0587_),
    .B2(_3226_),
    .Y(_2184_));
 sky130_fd_sc_hd__a221oi_1 _5760_ (.A1(_0593_),
    .A2(_3217_),
    .B1(_0563_),
    .B2(_3220_),
    .C1(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__nand2_1 _5761_ (.A(_3240_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_2186_));
 sky130_fd_sc_hd__o21ai_1 _5762_ (.A1(_0767_),
    .A2(_3237_),
    .B1(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__a221oi_1 _5763_ (.A1(_0549_),
    .A2(_3231_),
    .B1(_0558_),
    .B2(_3234_),
    .C1(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hd__nand2_1 _5764_ (.A(_3255_),
    .B(_3096_),
    .Y(_2189_));
 sky130_fd_sc_hd__o21ai_1 _5765_ (.A1(_3269_),
    .A2(_3252_),
    .B1(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__a221oi_1 _5766_ (.A1(_3099_),
    .A2(_3246_),
    .B1(_0619_),
    .B2(_3249_),
    .C1(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__o22ai_1 _5767_ (.A1(_0581_),
    .A2(_3267_),
    .B1(_0772_),
    .B2(_3270_),
    .Y(_2192_));
 sky130_fd_sc_hd__a221oi_1 _5768_ (.A1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .A2(_3261_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .B2(_3264_),
    .C1(_2192_),
    .Y(_2193_));
 sky130_fd_sc_hd__and4_1 _5769_ (.A(_2185_),
    .B(_2188_),
    .C(_2191_),
    .D(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__o22ai_1 _5770_ (.A1(_3398_),
    .A2(_3287_),
    .B1(_0690_),
    .B2(_3290_),
    .Y(_2195_));
 sky130_fd_sc_hd__a221oi_1 _5771_ (.A1(_0688_),
    .A2(_3280_),
    .B1(_3362_),
    .B2(_3284_),
    .C1(_2195_),
    .Y(_2196_));
 sky130_fd_sc_hd__nand2_1 _5772_ (.A(_3295_),
    .B(_3326_),
    .Y(_2197_));
 sky130_fd_sc_hd__nand2_1 _5773_ (.A(_3299_),
    .B(_3366_),
    .Y(_2198_));
 sky130_fd_sc_hd__nand2_1 _5774_ (.A(_3304_),
    .B(_0819_),
    .Y(_2199_));
 sky130_fd_sc_hd__nand2_1 _5775_ (.A(_3308_),
    .B(_3330_),
    .Y(_2200_));
 sky130_fd_sc_hd__and4_1 _5776_ (.A(_2197_),
    .B(_2198_),
    .C(_2199_),
    .D(_2200_),
    .X(_2201_));
 sky130_fd_sc_hd__o22ai_1 _5777_ (.A1(_1105_),
    .A2(_3313_),
    .B1(_1232_),
    .B2(_3316_),
    .Y(_2202_));
 sky130_fd_sc_hd__a22o_1 _5778_ (.A1(_3319_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .B1(_3321_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_2203_));
 sky130_fd_sc_hd__nor2_1 _5779_ (.A(_2202_),
    .B(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__o22ai_1 _5780_ (.A1(_0846_),
    .A2(_3335_),
    .B1(_0987_),
    .B2(_3338_),
    .Y(_2205_));
 sky130_fd_sc_hd__a221oi_1 _5781_ (.A1(_3350_),
    .A2(_3328_),
    .B1(_3403_),
    .B2(_3332_),
    .C1(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__and4_1 _5782_ (.A(_2196_),
    .B(_2201_),
    .C(_2204_),
    .D(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__nand2_1 _5783_ (.A(_3355_),
    .B(_3071_),
    .Y(_2208_));
 sky130_fd_sc_hd__nand2_1 _5784_ (.A(_3360_),
    .B(_3068_),
    .Y(_2209_));
 sky130_fd_sc_hd__nand2_1 _5785_ (.A(_2208_),
    .B(_2209_),
    .Y(_2210_));
 sky130_fd_sc_hd__a221oi_1 _5786_ (.A1(_3074_),
    .A2(_3348_),
    .B1(_3078_),
    .B2(_3352_),
    .C1(_2210_),
    .Y(_2211_));
 sky130_fd_sc_hd__nand2_1 _5787_ (.A(_3374_),
    .B(_3044_),
    .Y(_2212_));
 sky130_fd_sc_hd__nand2_1 _5788_ (.A(_3379_),
    .B(_0851_),
    .Y(_2213_));
 sky130_fd_sc_hd__nand2_1 _5789_ (.A(_2212_),
    .B(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__a221oi_1 _5790_ (.A1(_3407_),
    .A2(_3368_),
    .B1(_0693_),
    .B2(_3371_),
    .C1(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__nand2_1 _5791_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_2216_));
 sky130_fd_sc_hd__nand2_1 _5792_ (.A(_3394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_2217_));
 sky130_fd_sc_hd__or2_1 _5793_ (.A(_0811_),
    .B(_3399_),
    .X(_2218_));
 sky130_fd_sc_hd__o2111a_1 _5794_ (.A1(_3222_),
    .A2(_3386_),
    .B1(_2216_),
    .C1(_2217_),
    .D1(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__nand2_1 _5795_ (.A(_3415_),
    .B(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_2220_));
 sky130_fd_sc_hd__o21ai_1 _5796_ (.A1(_3266_),
    .A2(_3412_),
    .B1(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hd__a221oi_1 _5797_ (.A1(_3081_),
    .A2(_3405_),
    .B1(_3084_),
    .B2(_3409_),
    .C1(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__and4_1 _5798_ (.A(_2211_),
    .B(_2215_),
    .C(_2219_),
    .D(_2222_),
    .X(_2223_));
 sky130_fd_sc_hd__and4_1 _5799_ (.A(_2183_),
    .B(_2194_),
    .C(_2207_),
    .D(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(_0337_),
    .B(_0876_),
    .Y(_2225_));
 sky130_fd_sc_hd__nand2_1 _5801_ (.A(_0342_),
    .B(_0722_),
    .Y(_2226_));
 sky130_fd_sc_hd__nand2_1 _5802_ (.A(_2225_),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a221oi_1 _5803_ (.A1(_0720_),
    .A2(_0330_),
    .B1(_0874_),
    .B2(_0334_),
    .C1(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__o22ai_1 _5804_ (.A1(_0734_),
    .A2(_0349_),
    .B1(_0885_),
    .B2(_0352_),
    .Y(_2229_));
 sky130_fd_sc_hd__a22o_1 _5805_ (.A1(_0355_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .B1(_0358_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_2230_));
 sky130_fd_sc_hd__nor2_1 _5806_ (.A(_2229_),
    .B(_2230_),
    .Y(_2231_));
 sky130_fd_sc_hd__nand2_1 _5807_ (.A(_0375_),
    .B(_0869_),
    .Y(_2232_));
 sky130_fd_sc_hd__o21ai_1 _5808_ (.A1(_0389_),
    .A2(_0372_),
    .B1(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__a221oi_1 _5809_ (.A1(_0385_),
    .A2(_0365_),
    .B1(_0713_),
    .B2(_0369_),
    .C1(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(_0393_),
    .B(_0729_),
    .Y(_2235_));
 sky130_fd_sc_hd__o21ai_1 _5811_ (.A1(_0727_),
    .A2(_0390_),
    .B1(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__a221oi_1 _5812_ (.A1(_1012_),
    .A2(_0383_),
    .B1(_0427_),
    .B2(_0387_),
    .C1(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__and4_1 _5813_ (.A(_2228_),
    .B(_2231_),
    .C(_2234_),
    .D(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__nand2_1 _5814_ (.A(_0404_),
    .B(_3148_),
    .Y(_2239_));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(_0408_),
    .B(_3161_),
    .Y(_2240_));
 sky130_fd_sc_hd__or2_1 _5816_ (.A(_1070_),
    .B(_0413_),
    .X(_2241_));
 sky130_fd_sc_hd__o2111a_1 _5817_ (.A1(_0790_),
    .A2(_0401_),
    .B1(_2239_),
    .C1(_2240_),
    .D1(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__nand2_1 _5818_ (.A(_0421_),
    .B(_0630_),
    .Y(_2243_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_0425_),
    .B(_0632_),
    .Y(_2244_));
 sky130_fd_sc_hd__or2_1 _5820_ (.A(_0634_),
    .B(_0430_),
    .X(_2245_));
 sky130_fd_sc_hd__o2111a_1 _5821_ (.A1(_3123_),
    .A2(_0418_),
    .B1(_2243_),
    .C1(_2244_),
    .D1(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__nand2_1 _5822_ (.A(_0446_),
    .B(_0738_),
    .Y(_2247_));
 sky130_fd_sc_hd__o21ai_1 _5823_ (.A1(_0880_),
    .A2(_0443_),
    .B1(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__a221oi_1 _5824_ (.A1(_0889_),
    .A2(_0436_),
    .B1(_0890_),
    .B2(_0440_),
    .C1(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_0464_),
    .B(_3116_),
    .Y(_2250_));
 sky130_fd_sc_hd__o21ai_1 _5826_ (.A1(_0934_),
    .A2(_0461_),
    .B1(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__a221oi_1 _5827_ (.A1(_3131_),
    .A2(_0454_),
    .B1(_3104_),
    .B2(_0458_),
    .C1(_2251_),
    .Y(_2252_));
 sky130_fd_sc_hd__and4_1 _5828_ (.A(_2242_),
    .B(_2246_),
    .C(_2249_),
    .D(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__and2_1 _5829_ (.A(_2238_),
    .B(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__nand2_1 _5830_ (.A(_0478_),
    .B(_0357_),
    .Y(_2255_));
 sky130_fd_sc_hd__a22o_1 _5831_ (.A1(_0482_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .B1(_0484_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_2256_));
 sky130_fd_sc_hd__inv_2 _5832_ (.A(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__o211a_1 _5833_ (.A1(_0351_),
    .A2(_0475_),
    .B1(_2255_),
    .C1(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__nand2_1 _5834_ (.A(_0502_),
    .B(_0363_),
    .Y(_2259_));
 sky130_fd_sc_hd__o21ai_1 _5835_ (.A1(_1533_),
    .A2(_0499_),
    .B1(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__a221oi_1 _5836_ (.A1(_0539_),
    .A2(_0491_),
    .B1(_0528_),
    .B2(_0495_),
    .C1(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_0513_),
    .B(_0377_),
    .Y(_2262_));
 sky130_fd_sc_hd__nand2_1 _5838_ (.A(_0518_),
    .B(_0367_),
    .Y(_2263_));
 sky130_fd_sc_hd__or2_1 _5839_ (.A(_0371_),
    .B(_0524_),
    .X(_2264_));
 sky130_fd_sc_hd__o2111a_1 _5840_ (.A1(_0348_),
    .A2(_0510_),
    .B1(_2262_),
    .C1(_2263_),
    .D1(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__nand2_1 _5841_ (.A(_0537_),
    .B(_0326_),
    .Y(_2266_));
 sky130_fd_sc_hd__nand2_1 _5842_ (.A(_0542_),
    .B(_0339_),
    .Y(_2267_));
 sky130_fd_sc_hd__nand2_1 _5843_ (.A(_2266_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__a221oi_1 _5844_ (.A1(_0332_),
    .A2(_0530_),
    .B1(_0381_),
    .B2(_0534_),
    .C1(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__and4_1 _5845_ (.A(_2258_),
    .B(_2261_),
    .C(_2265_),
    .D(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(_0556_),
    .B(_0504_),
    .Y(_2271_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_0561_),
    .B(_0493_),
    .Y(_2272_));
 sky130_fd_sc_hd__or2_1 _5848_ (.A(_0901_),
    .B(_0566_),
    .X(_2273_));
 sky130_fd_sc_hd__o2111a_1 _5849_ (.A1(_0498_),
    .A2(_0553_),
    .B1(_2271_),
    .C1(_2272_),
    .D1(_2273_),
    .X(_2274_));
 sky130_fd_sc_hd__nand2_1 _5850_ (.A(_0574_),
    .B(_0508_),
    .Y(_2275_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_0578_),
    .B(_0522_),
    .Y(_2276_));
 sky130_fd_sc_hd__or2_1 _5852_ (.A(_0756_),
    .B(_0582_),
    .X(_2277_));
 sky130_fd_sc_hd__o2111a_1 _5853_ (.A1(_0472_),
    .A2(_0571_),
    .B1(_2275_),
    .C1(_2276_),
    .D1(_2277_),
    .X(_2278_));
 sky130_fd_sc_hd__or2_1 _5854_ (.A(_1058_),
    .B(_0595_),
    .X(_2279_));
 sky130_fd_sc_hd__o221a_1 _5855_ (.A1(_0924_),
    .A2(_0588_),
    .B1(_0778_),
    .B2(_0591_),
    .C1(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__o22ai_1 _5856_ (.A1(_0744_),
    .A2(_0606_),
    .B1(_0896_),
    .B2(_0609_),
    .Y(_2281_));
 sky130_fd_sc_hd__a221oi_1 _5857_ (.A1(_0486_),
    .A2(_0600_),
    .B1(_0544_),
    .B2(_0603_),
    .C1(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__and4_1 _5858_ (.A(_2274_),
    .B(_2278_),
    .C(_2280_),
    .D(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__and3_1 _5859_ (.A(_2254_),
    .B(_2270_),
    .C(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__nand2_1 _5860_ (.A(_0617_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_2285_));
 sky130_fd_sc_hd__nand3_1 _5861_ (.A(_2224_),
    .B(_2284_),
    .C(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__inv_2 _5862_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2287_));
 sky130_fd_sc_hd__a21oi_1 _5863_ (.A1(_2287_),
    .A2(_3102_),
    .B1(_2984_),
    .Y(_2288_));
 sky130_fd_sc_hd__o21a_1 _5864_ (.A1(_0932_),
    .A2(_2286_),
    .B1(_2288_),
    .X(_0284_));
 sky130_fd_sc_hd__o22ai_1 _5865_ (.A1(_0668_),
    .A2(_3129_),
    .B1(_0829_),
    .B2(_3137_),
    .Y(_2289_));
 sky130_fd_sc_hd__a221oi_1 _5866_ (.A1(_0670_),
    .A2(_3114_),
    .B1(_0831_),
    .B2(_3121_),
    .C1(_2289_),
    .Y(_2290_));
 sky130_fd_sc_hd__nand2_1 _5867_ (.A(_3159_),
    .B(_3195_),
    .Y(_2291_));
 sky130_fd_sc_hd__o21ai_1 _5868_ (.A1(_1195_),
    .A2(_3155_),
    .B1(_2291_),
    .Y(_2292_));
 sky130_fd_sc_hd__a221oi_1 _5869_ (.A1(_0637_),
    .A2(_3146_),
    .B1(_0799_),
    .B2(_3151_),
    .C1(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__nand2_1 _5870_ (.A(_3173_),
    .B(_0661_),
    .Y(_2294_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(_3179_),
    .B(_0663_),
    .Y(_2295_));
 sky130_fd_sc_hd__or2_1 _5872_ (.A(_1812_),
    .B(_3186_),
    .X(_2296_));
 sky130_fd_sc_hd__o2111a_1 _5873_ (.A1(_3315_),
    .A2(_3168_),
    .B1(_2294_),
    .C1(_2295_),
    .D1(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__nand2_1 _5874_ (.A(_3201_),
    .B(_3282_),
    .Y(_2298_));
 sky130_fd_sc_hd__nand2_1 _5875_ (.A(_3207_),
    .B(_3275_),
    .Y(_2299_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_2298_),
    .B(_2299_),
    .Y(_2300_));
 sky130_fd_sc_hd__a221oi_1 _5877_ (.A1(_0657_),
    .A2(_3193_),
    .B1(_0819_),
    .B2(_3197_),
    .C1(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__and4_1 _5878_ (.A(_2290_),
    .B(_2293_),
    .C(_2297_),
    .D(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__o22ai_1 _5879_ (.A1(_0587_),
    .A2(_3223_),
    .B1(_0594_),
    .B2(_3226_),
    .Y(_2303_));
 sky130_fd_sc_hd__a221oi_1 _5880_ (.A1(_0563_),
    .A2(_3217_),
    .B1(_0549_),
    .B2(_3220_),
    .C1(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__nand2_1 _5881_ (.A(_3240_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_2305_));
 sky130_fd_sc_hd__o21ai_1 _5882_ (.A1(_0581_),
    .A2(_3237_),
    .B1(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__a221oi_1 _5883_ (.A1(_0558_),
    .A2(_3231_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .B2(_3234_),
    .C1(_2306_),
    .Y(_2307_));
 sky130_fd_sc_hd__nand2_1 _5884_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_2308_));
 sky130_fd_sc_hd__o21ai_1 _5885_ (.A1(_0653_),
    .A2(_3252_),
    .B1(_2308_),
    .Y(_2309_));
 sky130_fd_sc_hd__a221oi_1 _5886_ (.A1(_0619_),
    .A2(_3246_),
    .B1(_0783_),
    .B2(_3249_),
    .C1(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__o22ai_1 _5887_ (.A1(_0772_),
    .A2(_3267_),
    .B1(_0570_),
    .B2(_3270_),
    .Y(_2311_));
 sky130_fd_sc_hd__a221oi_1 _5888_ (.A1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .A2(_3261_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .B2(_3264_),
    .C1(_2311_),
    .Y(_2312_));
 sky130_fd_sc_hd__and4_1 _5889_ (.A(_2304_),
    .B(_2307_),
    .C(_2310_),
    .D(_2312_),
    .X(_2313_));
 sky130_fd_sc_hd__o22ai_1 _5890_ (.A1(_0690_),
    .A2(_3287_),
    .B1(_3385_),
    .B2(_3290_),
    .Y(_2314_));
 sky130_fd_sc_hd__a221oi_1 _5891_ (.A1(_3362_),
    .A2(_3280_),
    .B1(_3357_),
    .B2(_3284_),
    .C1(_2314_),
    .Y(_2315_));
 sky130_fd_sc_hd__nand2_1 _5892_ (.A(_3295_),
    .B(_3330_),
    .Y(_2316_));
 sky130_fd_sc_hd__nand2_1 _5893_ (.A(_3299_),
    .B(_3370_),
    .Y(_2317_));
 sky130_fd_sc_hd__nand2_1 _5894_ (.A(_3304_),
    .B(_3326_),
    .Y(_2318_));
 sky130_fd_sc_hd__nand2_1 _5895_ (.A(_3308_),
    .B(_3366_),
    .Y(_2319_));
 sky130_fd_sc_hd__and4_1 _5896_ (.A(_2316_),
    .B(_2317_),
    .C(_2318_),
    .D(_2319_),
    .X(_2320_));
 sky130_fd_sc_hd__o22ai_1 _5897_ (.A1(_1232_),
    .A2(_3313_),
    .B1(_1356_),
    .B2(_3316_),
    .Y(_2321_));
 sky130_fd_sc_hd__a22o_1 _5898_ (.A1(_3319_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .B1(_3321_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_2322_));
 sky130_fd_sc_hd__nor2_1 _5899_ (.A(_2321_),
    .B(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__o22ai_1 _5900_ (.A1(_0987_),
    .A2(_3335_),
    .B1(_1117_),
    .B2(_3338_),
    .Y(_2324_));
 sky130_fd_sc_hd__a221oi_1 _5901_ (.A1(_3403_),
    .A2(_3328_),
    .B1(_3407_),
    .B2(_3332_),
    .C1(_2324_),
    .Y(_2325_));
 sky130_fd_sc_hd__and4_1 _5902_ (.A(_2315_),
    .B(_2320_),
    .C(_2323_),
    .D(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__nand2_1 _5903_ (.A(_3355_),
    .B(_3074_),
    .Y(_2327_));
 sky130_fd_sc_hd__nand2_1 _5904_ (.A(_3360_),
    .B(_3071_),
    .Y(_2328_));
 sky130_fd_sc_hd__nand2_1 _5905_ (.A(_2327_),
    .B(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__a221oi_1 _5906_ (.A1(_3078_),
    .A2(_3348_),
    .B1(_3081_),
    .B2(_3352_),
    .C1(_2329_),
    .Y(_2330_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(_3374_),
    .B(_3056_),
    .Y(_2331_));
 sky130_fd_sc_hd__nand2_1 _5908_ (.A(_3379_),
    .B(_3044_),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _5909_ (.A(_2331_),
    .B(_2332_),
    .Y(_2333_));
 sky130_fd_sc_hd__a221oi_1 _5910_ (.A1(_0693_),
    .A2(_3368_),
    .B1(_0851_),
    .B2(_3371_),
    .C1(_2333_),
    .Y(_2334_));
 sky130_fd_sc_hd__nand2_1 _5911_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_2335_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(_3394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_2336_));
 sky130_fd_sc_hd__or2_1 _5913_ (.A(_0956_),
    .B(_3399_),
    .X(_2337_));
 sky130_fd_sc_hd__o2111a_1 _5914_ (.A1(_3225_),
    .A2(_3386_),
    .B1(_2335_),
    .C1(_2336_),
    .D1(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__nand2_1 _5915_ (.A(_3415_),
    .B(_3090_),
    .Y(_2339_));
 sky130_fd_sc_hd__o21ai_1 _5916_ (.A1(_3269_),
    .A2(_3412_),
    .B1(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__a221oi_1 _5917_ (.A1(_3084_),
    .A2(_3405_),
    .B1(_3087_),
    .B2(_3409_),
    .C1(_2340_),
    .Y(_2341_));
 sky130_fd_sc_hd__and4_1 _5918_ (.A(_2330_),
    .B(_2334_),
    .C(_2338_),
    .D(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__and4_1 _5919_ (.A(_2302_),
    .B(_2313_),
    .C(_2326_),
    .D(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__nand2_1 _5920_ (.A(_0337_),
    .B(_0720_),
    .Y(_2344_));
 sky130_fd_sc_hd__nand2_1 _5921_ (.A(_0342_),
    .B(_0876_),
    .Y(_2345_));
 sky130_fd_sc_hd__nand2_1 _5922_ (.A(_2344_),
    .B(_2345_),
    .Y(_2346_));
 sky130_fd_sc_hd__a221oi_1 _5923_ (.A1(_0874_),
    .A2(_0330_),
    .B1(_1012_),
    .B2(_0334_),
    .C1(_2346_),
    .Y(_2347_));
 sky130_fd_sc_hd__o22ai_1 _5924_ (.A1(_0885_),
    .A2(_0349_),
    .B1(_1022_),
    .B2(_0352_),
    .Y(_2348_));
 sky130_fd_sc_hd__a22o_1 _5925_ (.A1(_0355_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .B1(_0358_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .X(_2349_));
 sky130_fd_sc_hd__nor2_1 _5926_ (.A(_2348_),
    .B(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__nand2_1 _5927_ (.A(_0375_),
    .B(_0448_),
    .Y(_2351_));
 sky130_fd_sc_hd__o21ai_1 _5928_ (.A1(_0442_),
    .A2(_0372_),
    .B1(_2351_),
    .Y(_2352_));
 sky130_fd_sc_hd__a221oi_1 _5929_ (.A1(_0713_),
    .A2(_0365_),
    .B1(_0714_),
    .B2(_0369_),
    .C1(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__nand2_1 _5930_ (.A(_0393_),
    .B(_0452_),
    .Y(_2354_));
 sky130_fd_sc_hd__o21ai_1 _5931_ (.A1(_0880_),
    .A2(_0390_),
    .B1(_2354_),
    .Y(_2355_));
 sky130_fd_sc_hd__a221oi_1 _5932_ (.A1(_0427_),
    .A2(_0383_),
    .B1(_0729_),
    .B2(_0387_),
    .C1(_2355_),
    .Y(_2356_));
 sky130_fd_sc_hd__and4_1 _5933_ (.A(_2347_),
    .B(_2350_),
    .C(_2353_),
    .D(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(_0404_),
    .B(_3175_),
    .Y(_2358_));
 sky130_fd_sc_hd__nand2_1 _5935_ (.A(_0408_),
    .B(_3141_),
    .Y(_2359_));
 sky130_fd_sc_hd__or2_1 _5936_ (.A(_3183_),
    .B(_0413_),
    .X(_2360_));
 sky130_fd_sc_hd__o2111a_1 _5937_ (.A1(_0937_),
    .A2(_0401_),
    .B1(_2358_),
    .C1(_2359_),
    .D1(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__nand2_1 _5938_ (.A(_0421_),
    .B(_3181_),
    .Y(_2362_));
 sky130_fd_sc_hd__nand2_1 _5939_ (.A(_0425_),
    .B(_0795_),
    .Y(_2363_));
 sky130_fd_sc_hd__or2_1 _5940_ (.A(_3165_),
    .B(_0430_),
    .X(_2364_));
 sky130_fd_sc_hd__o2111a_1 _5941_ (.A1(_3132_),
    .A2(_0418_),
    .B1(_2362_),
    .C1(_2363_),
    .D1(_2364_),
    .X(_2365_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_0446_),
    .B(_0889_),
    .Y(_2366_));
 sky130_fd_sc_hd__o21ai_1 _5943_ (.A1(_1017_),
    .A2(_0443_),
    .B1(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__a221oi_1 _5944_ (.A1(_0890_),
    .A2(_0436_),
    .B1(_3161_),
    .B2(_0440_),
    .C1(_2367_),
    .Y(_2368_));
 sky130_fd_sc_hd__nand2_1 _5945_ (.A(_0464_),
    .B(_3209_),
    .Y(_2369_));
 sky130_fd_sc_hd__o21ai_1 _5946_ (.A1(_1067_),
    .A2(_0461_),
    .B1(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__a221oi_1 _5947_ (.A1(_3104_),
    .A2(_0454_),
    .B1(_3116_),
    .B2(_0458_),
    .C1(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__and4_1 _5948_ (.A(_2361_),
    .B(_2365_),
    .C(_2368_),
    .D(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__and2_1 _5949_ (.A(_2357_),
    .B(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_0478_),
    .B(_0360_),
    .Y(_2374_));
 sky130_fd_sc_hd__a22o_1 _5951_ (.A1(_0482_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .B1(_0484_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_2375_));
 sky130_fd_sc_hd__inv_2 _5952_ (.A(_2375_),
    .Y(_2376_));
 sky130_fd_sc_hd__o211a_1 _5953_ (.A1(_0703_),
    .A2(_0475_),
    .B1(_2374_),
    .C1(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__nand2_1 _5954_ (.A(_0502_),
    .B(_0367_),
    .Y(_2378_));
 sky130_fd_sc_hd__o21ai_1 _5955_ (.A1(_1655_),
    .A2(_0499_),
    .B1(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__a221oi_1 _5956_ (.A1(_0528_),
    .A2(_0491_),
    .B1(_0532_),
    .B2(_0495_),
    .C1(_2379_),
    .Y(_2380_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(_0513_),
    .B(_0709_),
    .Y(_2381_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_0518_),
    .B(_0707_),
    .Y(_2382_));
 sky130_fd_sc_hd__or2_1 _5959_ (.A(_0708_),
    .B(_0524_),
    .X(_2383_));
 sky130_fd_sc_hd__o2111a_1 _5960_ (.A1(_0351_),
    .A2(_0510_),
    .B1(_2381_),
    .C1(_2382_),
    .D1(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__nand2_1 _5961_ (.A(_0537_),
    .B(_0332_),
    .Y(_2385_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(_0542_),
    .B(_0326_),
    .Y(_2386_));
 sky130_fd_sc_hd__nand2_1 _5963_ (.A(_2385_),
    .B(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__a221oi_1 _5964_ (.A1(_0381_),
    .A2(_0530_),
    .B1(_0385_),
    .B2(_0534_),
    .C1(_2387_),
    .Y(_2388_));
 sky130_fd_sc_hd__and4_1 _5965_ (.A(_2377_),
    .B(_2380_),
    .C(_2384_),
    .D(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__nand2_1 _5966_ (.A(_0556_),
    .B(_0520_),
    .Y(_2390_));
 sky130_fd_sc_hd__nand2_1 _5967_ (.A(_0561_),
    .B(_0497_),
    .Y(_2391_));
 sky130_fd_sc_hd__or2_1 _5968_ (.A(_0523_),
    .B(_0566_),
    .X(_2392_));
 sky130_fd_sc_hd__o2111a_1 _5969_ (.A1(_0750_),
    .A2(_0553_),
    .B1(_2390_),
    .C1(_2391_),
    .D1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__nand2_1 _5970_ (.A(_0574_),
    .B(_0471_),
    .Y(_2394_));
 sky130_fd_sc_hd__nand2_1 _5971_ (.A(_0578_),
    .B(_0515_),
    .Y(_2395_));
 sky130_fd_sc_hd__or2_1 _5972_ (.A(_0509_),
    .B(_0582_),
    .X(_2396_));
 sky130_fd_sc_hd__o2111a_1 _5973_ (.A1(_0744_),
    .A2(_0571_),
    .B1(_2394_),
    .C1(_2395_),
    .D1(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__or2_1 _5974_ (.A(_1186_),
    .B(_0595_),
    .X(_2398_));
 sky130_fd_sc_hd__o221a_1 _5975_ (.A1(_1058_),
    .A2(_0588_),
    .B1(_0924_),
    .B2(_0591_),
    .C1(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__o22ai_1 _5976_ (.A1(_0896_),
    .A2(_0606_),
    .B1(_1031_),
    .B2(_0609_),
    .Y(_2400_));
 sky130_fd_sc_hd__a221oi_1 _5977_ (.A1(_0544_),
    .A2(_0600_),
    .B1(_0539_),
    .B2(_0603_),
    .C1(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__and4_1 _5978_ (.A(_2393_),
    .B(_2397_),
    .C(_2399_),
    .D(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__and3_1 _5979_ (.A(_2373_),
    .B(_2389_),
    .C(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__nand2_1 _5980_ (.A(_0617_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_2404_));
 sky130_fd_sc_hd__nand3_1 _5981_ (.A(_2343_),
    .B(_2403_),
    .C(_2404_),
    .Y(_2405_));
 sky130_fd_sc_hd__inv_2 _5982_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2406_));
 sky130_fd_sc_hd__a21oi_1 _5983_ (.A1(_2406_),
    .A2(_3102_),
    .B1(_2984_),
    .Y(_2407_));
 sky130_fd_sc_hd__o21a_1 _5984_ (.A1(_0932_),
    .A2(_2405_),
    .B1(_2407_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(_3050_),
    .B(_3024_),
    .Y(_2408_));
 sky130_fd_sc_hd__and3_1 _5986_ (.A(_3053_),
    .B(_3035_),
    .C(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__clkbuf_1 _5987_ (.A(_2409_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _5988_ (.A(_3049_),
    .B(_3017_),
    .Y(_2410_));
 sky130_fd_sc_hd__and3_1 _5989_ (.A(_3050_),
    .B(_3035_),
    .C(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__clkbuf_1 _5990_ (.A(_2411_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _5991_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .B(_3048_),
    .X(_2412_));
 sky130_fd_sc_hd__and3_1 _5992_ (.A(_2412_),
    .B(_3035_),
    .C(_3049_),
    .X(_2413_));
 sky130_fd_sc_hd__clkbuf_1 _5993_ (.A(_2413_),
    .X(_0280_));
 sky130_fd_sc_hd__nand2_4 _5994_ (.A(_3048_),
    .B(_3025_),
    .Y(_2414_));
 sky130_fd_sc_hd__clkbuf_4 _5995_ (.A(_2414_),
    .X(_2415_));
 sky130_fd_sc_hd__mux2_1 _5996_ (.A0(net7),
    .A1(_0619_),
    .S(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__and2_1 _5997_ (.A(_2416_),
    .B(_3076_),
    .X(_2417_));
 sky130_fd_sc_hd__clkbuf_1 _5998_ (.A(_2417_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5999_ (.A0(net6),
    .A1(_0783_),
    .S(_2415_),
    .X(_2418_));
 sky130_fd_sc_hd__clkbuf_2 _6000_ (.A(_3035_),
    .X(_2419_));
 sky130_fd_sc_hd__and2_1 _6001_ (.A(_2418_),
    .B(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__clkbuf_1 _6002_ (.A(_2420_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _6003_ (.A0(net5),
    .A1(_0586_),
    .S(_2415_),
    .X(_2421_));
 sky130_fd_sc_hd__and2_1 _6004_ (.A(_2421_),
    .B(_2419_),
    .X(_2422_));
 sky130_fd_sc_hd__clkbuf_1 _6005_ (.A(_2422_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _6006_ (.A0(net4),
    .A1(_0593_),
    .S(_2415_),
    .X(_2423_));
 sky130_fd_sc_hd__and2_1 _6007_ (.A(_2423_),
    .B(_2419_),
    .X(_2424_));
 sky130_fd_sc_hd__clkbuf_1 _6008_ (.A(_2424_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _6009_ (.A0(net3),
    .A1(_0563_),
    .S(_2415_),
    .X(_2425_));
 sky130_fd_sc_hd__and2_1 _6010_ (.A(_2425_),
    .B(_2419_),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _6011_ (.A(_2426_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _6012_ (.A0(net2),
    .A1(_0549_),
    .S(_2415_),
    .X(_2427_));
 sky130_fd_sc_hd__and2_1 _6013_ (.A(_2427_),
    .B(_2419_),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_1 _6014_ (.A(_2428_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _6015_ (.A0(net16),
    .A1(_0558_),
    .S(_2415_),
    .X(_2429_));
 sky130_fd_sc_hd__and2_1 _6016_ (.A(_2429_),
    .B(_2419_),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_1 _6017_ (.A(_2430_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _6018_ (.A0(net15),
    .A1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .S(_2415_),
    .X(_2431_));
 sky130_fd_sc_hd__and2_1 _6019_ (.A(_2431_),
    .B(_2419_),
    .X(_2432_));
 sky130_fd_sc_hd__clkbuf_1 _6020_ (.A(_2432_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _6021_ (.A0(net14),
    .A1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .S(_2415_),
    .X(_2433_));
 sky130_fd_sc_hd__and2_1 _6022_ (.A(_2433_),
    .B(_2419_),
    .X(_2434_));
 sky130_fd_sc_hd__clkbuf_1 _6023_ (.A(_2434_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _6024_ (.A0(net13),
    .A1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .S(_2415_),
    .X(_2435_));
 sky130_fd_sc_hd__and2_1 _6025_ (.A(_2435_),
    .B(_2419_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_1 _6026_ (.A(_2436_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _6027_ (.A0(net12),
    .A1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .S(_2414_),
    .X(_2437_));
 sky130_fd_sc_hd__and2_1 _6028_ (.A(_2437_),
    .B(_2419_),
    .X(_2438_));
 sky130_fd_sc_hd__clkbuf_1 _6029_ (.A(_2438_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _6030_ (.A0(net11),
    .A1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .S(_2414_),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_2 _6031_ (.A(_3035_),
    .X(_2440_));
 sky130_fd_sc_hd__and2_1 _6032_ (.A(_2439_),
    .B(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__clkbuf_1 _6033_ (.A(_2441_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(net10),
    .A1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .S(_2414_),
    .X(_2442_));
 sky130_fd_sc_hd__and2_1 _6035_ (.A(_2442_),
    .B(_2440_),
    .X(_2443_));
 sky130_fd_sc_hd__clkbuf_1 _6036_ (.A(_2443_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _6037_ (.A0(net9),
    .A1(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .S(_2414_),
    .X(_2444_));
 sky130_fd_sc_hd__and2_1 _6038_ (.A(_2444_),
    .B(_2440_),
    .X(_2445_));
 sky130_fd_sc_hd__clkbuf_1 _6039_ (.A(_2445_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _6040_ (.A0(net8),
    .A1(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .S(_2414_),
    .X(_2446_));
 sky130_fd_sc_hd__and2_1 _6041_ (.A(_2446_),
    .B(_2440_),
    .X(_2447_));
 sky130_fd_sc_hd__clkbuf_1 _6042_ (.A(_2447_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _6043_ (.A0(net1),
    .A1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .S(_2414_),
    .X(_2448_));
 sky130_fd_sc_hd__and2_1 _6044_ (.A(_2448_),
    .B(_2440_),
    .X(_2449_));
 sky130_fd_sc_hd__clkbuf_1 _6045_ (.A(_2449_),
    .X(_0264_));
 sky130_fd_sc_hd__or4b_1 _6046_ (.A(net196),
    .B(net198),
    .C(_3018_),
    .D_N(_3048_),
    .X(_2450_));
 sky130_fd_sc_hd__buf_2 _6047_ (.A(net199),
    .X(_2451_));
 sky130_fd_sc_hd__clkbuf_4 _6048_ (.A(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_1 _6049_ (.A0(net7),
    .A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .S(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__and2_1 _6050_ (.A(_2453_),
    .B(_2440_),
    .X(_2454_));
 sky130_fd_sc_hd__clkbuf_1 _6051_ (.A(_2454_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _6052_ (.A0(net6),
    .A1(_0493_),
    .S(_2452_),
    .X(_2455_));
 sky130_fd_sc_hd__and2_1 _6053_ (.A(_2455_),
    .B(_2440_),
    .X(_2456_));
 sky130_fd_sc_hd__clkbuf_1 _6054_ (.A(_2456_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _6055_ (.A0(net5),
    .A1(_0497_),
    .S(_2452_),
    .X(_2457_));
 sky130_fd_sc_hd__and2_1 _6056_ (.A(_2457_),
    .B(_2440_),
    .X(_2458_));
 sky130_fd_sc_hd__clkbuf_1 _6057_ (.A(_2458_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _6058_ (.A0(net4),
    .A1(_0504_),
    .S(_2452_),
    .X(_2459_));
 sky130_fd_sc_hd__and2_1 _6059_ (.A(_2459_),
    .B(_2440_),
    .X(_2460_));
 sky130_fd_sc_hd__clkbuf_1 _6060_ (.A(_2460_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _6061_ (.A0(net3),
    .A1(_0520_),
    .S(_2452_),
    .X(_2461_));
 sky130_fd_sc_hd__and2_1 _6062_ (.A(_2461_),
    .B(_2440_),
    .X(_2462_));
 sky130_fd_sc_hd__clkbuf_1 _6063_ (.A(_2462_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _6064_ (.A0(net2),
    .A1(_0522_),
    .S(_2452_),
    .X(_2463_));
 sky130_fd_sc_hd__clkbuf_2 _6065_ (.A(_3035_),
    .X(_2464_));
 sky130_fd_sc_hd__and2_1 _6066_ (.A(_2463_),
    .B(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__clkbuf_1 _6067_ (.A(_2465_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _6068_ (.A0(net16),
    .A1(_0515_),
    .S(_2452_),
    .X(_2466_));
 sky130_fd_sc_hd__and2_1 _6069_ (.A(_2466_),
    .B(_2464_),
    .X(_2467_));
 sky130_fd_sc_hd__clkbuf_1 _6070_ (.A(_2467_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _6071_ (.A0(net15),
    .A1(_0508_),
    .S(_2452_),
    .X(_2468_));
 sky130_fd_sc_hd__and2_1 _6072_ (.A(_2468_),
    .B(_2464_),
    .X(_2469_));
 sky130_fd_sc_hd__clkbuf_1 _6073_ (.A(_2469_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _6074_ (.A0(net14),
    .A1(_0471_),
    .S(_2452_),
    .X(_2470_));
 sky130_fd_sc_hd__and2_1 _6075_ (.A(_2470_),
    .B(_2464_),
    .X(_2471_));
 sky130_fd_sc_hd__clkbuf_1 _6076_ (.A(_2471_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _6077_ (.A0(net13),
    .A1(_0480_),
    .S(_2452_),
    .X(_2472_));
 sky130_fd_sc_hd__and2_1 _6078_ (.A(_2472_),
    .B(_2464_),
    .X(_2473_));
 sky130_fd_sc_hd__clkbuf_1 _6079_ (.A(_2473_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _6080_ (.A0(net12),
    .A1(_0745_),
    .S(_2451_),
    .X(_2474_));
 sky130_fd_sc_hd__and2_1 _6081_ (.A(_2474_),
    .B(_2464_),
    .X(_2475_));
 sky130_fd_sc_hd__clkbuf_1 _6082_ (.A(_2475_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _6083_ (.A0(net11),
    .A1(_0486_),
    .S(_2451_),
    .X(_2476_));
 sky130_fd_sc_hd__and2_1 _6084_ (.A(_2476_),
    .B(_2464_),
    .X(_2477_));
 sky130_fd_sc_hd__clkbuf_1 _6085_ (.A(_2477_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _6086_ (.A0(net10),
    .A1(_0544_),
    .S(_2451_),
    .X(_2478_));
 sky130_fd_sc_hd__and2_1 _6087_ (.A(_2478_),
    .B(_2464_),
    .X(_2479_));
 sky130_fd_sc_hd__clkbuf_1 _6088_ (.A(_2479_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _6089_ (.A0(net9),
    .A1(_0539_),
    .S(_2451_),
    .X(_2480_));
 sky130_fd_sc_hd__and2_1 _6090_ (.A(_2480_),
    .B(_2464_),
    .X(_2481_));
 sky130_fd_sc_hd__clkbuf_1 _6091_ (.A(_2481_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _6092_ (.A0(net8),
    .A1(_0528_),
    .S(_2451_),
    .X(_2482_));
 sky130_fd_sc_hd__and2_1 _6093_ (.A(_2482_),
    .B(_2464_),
    .X(_2483_));
 sky130_fd_sc_hd__clkbuf_1 _6094_ (.A(_2483_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _6095_ (.A0(net1),
    .A1(_0532_),
    .S(_2451_),
    .X(_2484_));
 sky130_fd_sc_hd__buf_2 _6096_ (.A(_3035_),
    .X(_2485_));
 sky130_fd_sc_hd__and2_1 _6097_ (.A(_2484_),
    .B(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__clkbuf_1 _6098_ (.A(_2486_),
    .X(_0248_));
 sky130_fd_sc_hd__or4b_2 _6099_ (.A(net196),
    .B(_3017_),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .D_N(_3048_),
    .X(_2487_));
 sky130_fd_sc_hd__buf_2 _6100_ (.A(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__buf_4 _6101_ (.A(_2488_),
    .X(_2489_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(net7),
    .A1(_0363_),
    .S(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__and2_1 _6103_ (.A(_2490_),
    .B(_2485_),
    .X(_2491_));
 sky130_fd_sc_hd__clkbuf_1 _6104_ (.A(_2491_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _6105_ (.A0(net6),
    .A1(_0367_),
    .S(_2489_),
    .X(_2492_));
 sky130_fd_sc_hd__and2_1 _6106_ (.A(_2492_),
    .B(_2485_),
    .X(_2493_));
 sky130_fd_sc_hd__clkbuf_1 _6107_ (.A(_2493_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _6108_ (.A0(net5),
    .A1(_0707_),
    .S(_2489_),
    .X(_2494_));
 sky130_fd_sc_hd__and2_1 _6109_ (.A(_2494_),
    .B(_2485_),
    .X(_2495_));
 sky130_fd_sc_hd__clkbuf_1 _6110_ (.A(_2495_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _6111_ (.A0(net4),
    .A1(_0377_),
    .S(_2489_),
    .X(_2496_));
 sky130_fd_sc_hd__and2_1 _6112_ (.A(_2496_),
    .B(_2485_),
    .X(_2497_));
 sky130_fd_sc_hd__clkbuf_1 _6113_ (.A(_2497_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _6114_ (.A0(net3),
    .A1(_0709_),
    .S(_2489_),
    .X(_2498_));
 sky130_fd_sc_hd__and2_1 _6115_ (.A(_2498_),
    .B(_2485_),
    .X(_2499_));
 sky130_fd_sc_hd__clkbuf_1 _6116_ (.A(_2499_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _6117_ (.A0(net2),
    .A1(_0865_),
    .S(_2489_),
    .X(_2500_));
 sky130_fd_sc_hd__and2_1 _6118_ (.A(_2500_),
    .B(_2485_),
    .X(_2501_));
 sky130_fd_sc_hd__clkbuf_1 _6119_ (.A(_2501_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _6120_ (.A0(net16),
    .A1(_0357_),
    .S(_2489_),
    .X(_2502_));
 sky130_fd_sc_hd__and2_1 _6121_ (.A(_2502_),
    .B(_2485_),
    .X(_2503_));
 sky130_fd_sc_hd__clkbuf_1 _6122_ (.A(_2503_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _6123_ (.A0(net15),
    .A1(_0360_),
    .S(_2489_),
    .X(_2504_));
 sky130_fd_sc_hd__and2_1 _6124_ (.A(_2504_),
    .B(_2485_),
    .X(_2505_));
 sky130_fd_sc_hd__clkbuf_1 _6125_ (.A(_2505_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _6126_ (.A0(net14),
    .A1(_0344_),
    .S(_2489_),
    .X(_2506_));
 sky130_fd_sc_hd__and2_1 _6127_ (.A(_2506_),
    .B(_2485_),
    .X(_2507_));
 sky130_fd_sc_hd__clkbuf_1 _6128_ (.A(_2507_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _6129_ (.A0(net13),
    .A1(_0339_),
    .S(_2489_),
    .X(_2508_));
 sky130_fd_sc_hd__clkbuf_2 _6130_ (.A(net19),
    .X(_2509_));
 sky130_fd_sc_hd__and2_1 _6131_ (.A(_2508_),
    .B(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__clkbuf_1 _6132_ (.A(_2510_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _6133_ (.A0(net12),
    .A1(_0326_),
    .S(_2488_),
    .X(_2511_));
 sky130_fd_sc_hd__and2_1 _6134_ (.A(_2511_),
    .B(_2509_),
    .X(_2512_));
 sky130_fd_sc_hd__clkbuf_1 _6135_ (.A(_2512_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _6136_ (.A0(net11),
    .A1(_0332_),
    .S(_2488_),
    .X(_2513_));
 sky130_fd_sc_hd__and2_1 _6137_ (.A(_2513_),
    .B(_2509_),
    .X(_2514_));
 sky130_fd_sc_hd__clkbuf_1 _6138_ (.A(_2514_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _6139_ (.A0(net10),
    .A1(_0381_),
    .S(_2488_),
    .X(_2515_));
 sky130_fd_sc_hd__and2_1 _6140_ (.A(_2515_),
    .B(_2509_),
    .X(_2516_));
 sky130_fd_sc_hd__clkbuf_1 _6141_ (.A(_2516_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _6142_ (.A0(net9),
    .A1(_0385_),
    .S(_2488_),
    .X(_2517_));
 sky130_fd_sc_hd__and2_1 _6143_ (.A(_2517_),
    .B(_2509_),
    .X(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _6144_ (.A(_2518_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _6145_ (.A0(net8),
    .A1(_0713_),
    .S(_2488_),
    .X(_2519_));
 sky130_fd_sc_hd__and2_1 _6146_ (.A(_2519_),
    .B(_2509_),
    .X(_2520_));
 sky130_fd_sc_hd__clkbuf_1 _6147_ (.A(_2520_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _6148_ (.A0(net1),
    .A1(_0714_),
    .S(_2488_),
    .X(_2521_));
 sky130_fd_sc_hd__and2_1 _6149_ (.A(_2521_),
    .B(_2509_),
    .X(_2522_));
 sky130_fd_sc_hd__clkbuf_1 _6150_ (.A(_2522_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_2 _6151_ (.A(net201),
    .B(_3050_),
    .X(_2523_));
 sky130_fd_sc_hd__buf_2 _6152_ (.A(_2523_),
    .X(_2524_));
 sky130_fd_sc_hd__clkbuf_4 _6153_ (.A(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__mux2_1 _6154_ (.A0(net7),
    .A1(_0869_),
    .S(_2525_),
    .X(_2526_));
 sky130_fd_sc_hd__and2_1 _6155_ (.A(_2526_),
    .B(_2509_),
    .X(_2527_));
 sky130_fd_sc_hd__clkbuf_1 _6156_ (.A(_2527_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _6157_ (.A0(net6),
    .A1(_0448_),
    .S(_2525_),
    .X(_2528_));
 sky130_fd_sc_hd__and2_1 _6158_ (.A(_2528_),
    .B(_2509_),
    .X(_2529_));
 sky130_fd_sc_hd__clkbuf_1 _6159_ (.A(_2529_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _6160_ (.A0(net5),
    .A1(_0434_),
    .S(_2525_),
    .X(_2530_));
 sky130_fd_sc_hd__and2_1 _6161_ (.A(_2530_),
    .B(_2509_),
    .X(_2531_));
 sky130_fd_sc_hd__clkbuf_1 _6162_ (.A(_2531_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _6163_ (.A0(net4),
    .A1(_0438_),
    .S(_2525_),
    .X(_2532_));
 sky130_fd_sc_hd__clkbuf_2 _6164_ (.A(net19),
    .X(_2533_));
 sky130_fd_sc_hd__and2_1 _6165_ (.A(_2532_),
    .B(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__clkbuf_1 _6166_ (.A(_2534_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _6167_ (.A0(net3),
    .A1(_0410_),
    .S(_2525_),
    .X(_2535_));
 sky130_fd_sc_hd__and2_1 _6168_ (.A(_2535_),
    .B(_2533_),
    .X(_2536_));
 sky130_fd_sc_hd__clkbuf_1 _6169_ (.A(_2536_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _6170_ (.A0(net2),
    .A1(_0722_),
    .S(_2525_),
    .X(_2537_));
 sky130_fd_sc_hd__and2_1 _6171_ (.A(_2537_),
    .B(_2533_),
    .X(_2538_));
 sky130_fd_sc_hd__clkbuf_1 _6172_ (.A(_2538_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _6173_ (.A0(net16),
    .A1(_0876_),
    .S(_2525_),
    .X(_2539_));
 sky130_fd_sc_hd__and2_1 _6174_ (.A(_2539_),
    .B(_2533_),
    .X(_2540_));
 sky130_fd_sc_hd__clkbuf_1 _6175_ (.A(_2540_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _6176_ (.A0(net15),
    .A1(_0720_),
    .S(_2525_),
    .X(_2541_));
 sky130_fd_sc_hd__and2_1 _6177_ (.A(_2541_),
    .B(_2533_),
    .X(_2542_));
 sky130_fd_sc_hd__clkbuf_1 _6178_ (.A(_2542_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _6179_ (.A0(net14),
    .A1(_0874_),
    .S(_2525_),
    .X(_2543_));
 sky130_fd_sc_hd__and2_1 _6180_ (.A(_2543_),
    .B(_2533_),
    .X(_2544_));
 sky130_fd_sc_hd__clkbuf_1 _6181_ (.A(_2544_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _6182_ (.A0(net13),
    .A1(_1012_),
    .S(_2525_),
    .X(_2545_));
 sky130_fd_sc_hd__and2_1 _6183_ (.A(_2545_),
    .B(_2533_),
    .X(_2546_));
 sky130_fd_sc_hd__clkbuf_1 _6184_ (.A(_2546_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _6185_ (.A0(net12),
    .A1(_0427_),
    .S(_2524_),
    .X(_2547_));
 sky130_fd_sc_hd__and2_1 _6186_ (.A(_2547_),
    .B(_2533_),
    .X(_2548_));
 sky130_fd_sc_hd__clkbuf_1 _6187_ (.A(_2548_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _6188_ (.A0(net11),
    .A1(_0729_),
    .S(_2524_),
    .X(_2549_));
 sky130_fd_sc_hd__and2_1 _6189_ (.A(_2549_),
    .B(_2533_),
    .X(_2550_));
 sky130_fd_sc_hd__clkbuf_1 _6190_ (.A(_2550_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _6191_ (.A0(net10),
    .A1(_0452_),
    .S(_2524_),
    .X(_2551_));
 sky130_fd_sc_hd__and2_1 _6192_ (.A(_2551_),
    .B(_2533_),
    .X(_2552_));
 sky130_fd_sc_hd__clkbuf_1 _6193_ (.A(_2552_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _6194_ (.A0(net9),
    .A1(_0456_),
    .S(_2524_),
    .X(_2553_));
 sky130_fd_sc_hd__clkbuf_2 _6195_ (.A(net19),
    .X(_2554_));
 sky130_fd_sc_hd__and2_1 _6196_ (.A(_2553_),
    .B(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__clkbuf_1 _6197_ (.A(_2555_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _6198_ (.A0(net8),
    .A1(_0738_),
    .S(_2524_),
    .X(_2556_));
 sky130_fd_sc_hd__and2_1 _6199_ (.A(_2556_),
    .B(_2554_),
    .X(_2557_));
 sky130_fd_sc_hd__clkbuf_1 _6200_ (.A(_2557_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _6201_ (.A0(net1),
    .A1(_0889_),
    .S(_2524_),
    .X(_2558_));
 sky130_fd_sc_hd__and2_1 _6202_ (.A(_2558_),
    .B(_2554_),
    .X(_2559_));
 sky130_fd_sc_hd__clkbuf_1 _6203_ (.A(_2559_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_4 _6204_ (.A(_3048_),
    .B(net197),
    .Y(_2560_));
 sky130_fd_sc_hd__clkbuf_4 _6205_ (.A(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__mux2_1 _6206_ (.A0(net7),
    .A1(_0890_),
    .S(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__and2_1 _6207_ (.A(_2562_),
    .B(_2554_),
    .X(_2563_));
 sky130_fd_sc_hd__clkbuf_1 _6208_ (.A(_2563_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _6209_ (.A0(net6),
    .A1(_3161_),
    .S(_2561_),
    .X(_2564_));
 sky130_fd_sc_hd__and2_1 _6210_ (.A(_2564_),
    .B(_2554_),
    .X(_2565_));
 sky130_fd_sc_hd__clkbuf_1 _6211_ (.A(_2565_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _6212_ (.A0(net5),
    .A1(_3141_),
    .S(_2561_),
    .X(_2566_));
 sky130_fd_sc_hd__and2_1 _6213_ (.A(_2566_),
    .B(_2554_),
    .X(_2567_));
 sky130_fd_sc_hd__clkbuf_1 _6214_ (.A(_2567_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _6215_ (.A0(net4),
    .A1(_3148_),
    .S(_2561_),
    .X(_2568_));
 sky130_fd_sc_hd__and2_1 _6216_ (.A(_2568_),
    .B(_2554_),
    .X(_2569_));
 sky130_fd_sc_hd__clkbuf_1 _6217_ (.A(_2569_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _6218_ (.A0(net3),
    .A1(_3175_),
    .S(_2561_),
    .X(_2570_));
 sky130_fd_sc_hd__and2_1 _6219_ (.A(_2570_),
    .B(_2554_),
    .X(_2571_));
 sky130_fd_sc_hd__clkbuf_1 _6220_ (.A(_2571_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _6221_ (.A0(net2),
    .A1(_0630_),
    .S(_2561_),
    .X(_2572_));
 sky130_fd_sc_hd__and2_1 _6222_ (.A(_2572_),
    .B(_2554_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_1 _6223_ (.A(_2573_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _6224_ (.A0(net16),
    .A1(_3181_),
    .S(_2561_),
    .X(_2574_));
 sky130_fd_sc_hd__and2_1 _6225_ (.A(_2574_),
    .B(_2554_),
    .X(_2575_));
 sky130_fd_sc_hd__clkbuf_1 _6226_ (.A(_2575_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _6227_ (.A0(net15),
    .A1(_0632_),
    .S(_2561_),
    .X(_2576_));
 sky130_fd_sc_hd__buf_2 _6228_ (.A(net19),
    .X(_2577_));
 sky130_fd_sc_hd__and2_1 _6229_ (.A(_2576_),
    .B(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__clkbuf_1 _6230_ (.A(_2578_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _6231_ (.A0(net14),
    .A1(_0795_),
    .S(_2561_),
    .X(_2579_));
 sky130_fd_sc_hd__and2_1 _6232_ (.A(_2579_),
    .B(_2577_),
    .X(_2580_));
 sky130_fd_sc_hd__clkbuf_1 _6233_ (.A(_2580_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _6234_ (.A0(net13),
    .A1(_3131_),
    .S(_2561_),
    .X(_2581_));
 sky130_fd_sc_hd__and2_1 _6235_ (.A(_2581_),
    .B(_2577_),
    .X(_2582_));
 sky130_fd_sc_hd__clkbuf_1 _6236_ (.A(_2582_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _6237_ (.A0(net12),
    .A1(_3104_),
    .S(_2560_),
    .X(_2583_));
 sky130_fd_sc_hd__and2_1 _6238_ (.A(_2583_),
    .B(_2577_),
    .X(_2584_));
 sky130_fd_sc_hd__clkbuf_1 _6239_ (.A(_2584_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _6240_ (.A0(net11),
    .A1(_3116_),
    .S(_2560_),
    .X(_2585_));
 sky130_fd_sc_hd__and2_1 _6241_ (.A(_2585_),
    .B(_2577_),
    .X(_2586_));
 sky130_fd_sc_hd__clkbuf_1 _6242_ (.A(_2586_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _6243_ (.A0(net10),
    .A1(_3209_),
    .S(_2560_),
    .X(_2587_));
 sky130_fd_sc_hd__and2_1 _6244_ (.A(_2587_),
    .B(_2577_),
    .X(_2588_));
 sky130_fd_sc_hd__clkbuf_1 _6245_ (.A(_2588_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _6246_ (.A0(net9),
    .A1(_3203_),
    .S(_2560_),
    .X(_2589_));
 sky130_fd_sc_hd__and2_1 _6247_ (.A(_2589_),
    .B(_2577_),
    .X(_2590_));
 sky130_fd_sc_hd__clkbuf_1 _6248_ (.A(_2590_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _6249_ (.A0(net8),
    .A1(_3190_),
    .S(_2560_),
    .X(_2591_));
 sky130_fd_sc_hd__and2_1 _6250_ (.A(_2591_),
    .B(_2577_),
    .X(_2592_));
 sky130_fd_sc_hd__clkbuf_1 _6251_ (.A(_2592_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _6252_ (.A0(net1),
    .A1(_3195_),
    .S(_2560_),
    .X(_2593_));
 sky130_fd_sc_hd__and2_1 _6253_ (.A(_2593_),
    .B(_2577_),
    .X(_2594_));
 sky130_fd_sc_hd__clkbuf_1 _6254_ (.A(_2594_),
    .X(_0200_));
 sky130_fd_sc_hd__or4b_1 _6255_ (.A(_3024_),
    .B(_3017_),
    .C(net200),
    .D_N(_3048_),
    .X(_2595_));
 sky130_fd_sc_hd__buf_2 _6256_ (.A(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__clkbuf_4 _6257_ (.A(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__mux2_1 _6258_ (.A0(net7),
    .A1(_3366_),
    .S(_2597_),
    .X(_2598_));
 sky130_fd_sc_hd__and2_1 _6259_ (.A(_2598_),
    .B(_2577_),
    .X(_2599_));
 sky130_fd_sc_hd__clkbuf_1 _6260_ (.A(_2599_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _6261_ (.A0(net6),
    .A1(_3370_),
    .S(_2597_),
    .X(_2600_));
 sky130_fd_sc_hd__clkbuf_2 _6262_ (.A(net19),
    .X(_2601_));
 sky130_fd_sc_hd__and2_1 _6263_ (.A(_2600_),
    .B(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__clkbuf_1 _6264_ (.A(_2602_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _6265_ (.A0(net5),
    .A1(_3381_),
    .S(_2597_),
    .X(_2603_));
 sky130_fd_sc_hd__and2_1 _6266_ (.A(_2603_),
    .B(_2601_),
    .X(_2604_));
 sky130_fd_sc_hd__clkbuf_1 _6267_ (.A(_2604_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _6268_ (.A0(net4),
    .A1(_3376_),
    .S(_2597_),
    .X(_2605_));
 sky130_fd_sc_hd__and2_1 _6269_ (.A(_2605_),
    .B(_2601_),
    .X(_2606_));
 sky130_fd_sc_hd__clkbuf_1 _6270_ (.A(_2606_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _6271_ (.A0(net3),
    .A1(_3391_),
    .S(_2597_),
    .X(_2607_));
 sky130_fd_sc_hd__and2_1 _6272_ (.A(_2607_),
    .B(_2601_),
    .X(_2608_));
 sky130_fd_sc_hd__clkbuf_1 _6273_ (.A(_2608_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _6274_ (.A0(net2),
    .A1(_0686_),
    .S(_2597_),
    .X(_2609_));
 sky130_fd_sc_hd__and2_1 _6275_ (.A(_2609_),
    .B(_2601_),
    .X(_2610_));
 sky130_fd_sc_hd__clkbuf_1 _6276_ (.A(_2610_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _6277_ (.A0(net16),
    .A1(_3396_),
    .S(_2597_),
    .X(_2611_));
 sky130_fd_sc_hd__and2_1 _6278_ (.A(_2611_),
    .B(_2601_),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_1 _6279_ (.A(_2612_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _6280_ (.A0(net15),
    .A1(_0688_),
    .S(_2597_),
    .X(_2613_));
 sky130_fd_sc_hd__and2_1 _6281_ (.A(_2613_),
    .B(_2601_),
    .X(_2614_));
 sky130_fd_sc_hd__clkbuf_1 _6282_ (.A(_2614_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _6283_ (.A0(net14),
    .A1(_3362_),
    .S(_2597_),
    .X(_2615_));
 sky130_fd_sc_hd__and2_1 _6284_ (.A(_2615_),
    .B(_2601_),
    .X(_2616_));
 sky130_fd_sc_hd__clkbuf_1 _6285_ (.A(_2616_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _6286_ (.A0(net13),
    .A1(_3357_),
    .S(_2597_),
    .X(_2617_));
 sky130_fd_sc_hd__and2_1 _6287_ (.A(_2617_),
    .B(_2601_),
    .X(_2618_));
 sky130_fd_sc_hd__clkbuf_1 _6288_ (.A(_2618_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _6289_ (.A0(net12),
    .A1(_3343_),
    .S(_2596_),
    .X(_2619_));
 sky130_fd_sc_hd__and2_1 _6290_ (.A(_2619_),
    .B(_2601_),
    .X(_2620_));
 sky130_fd_sc_hd__clkbuf_1 _6291_ (.A(_2620_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _6292_ (.A0(net11),
    .A1(_3350_),
    .S(_2596_),
    .X(_2621_));
 sky130_fd_sc_hd__buf_2 _6293_ (.A(net19),
    .X(_2622_));
 sky130_fd_sc_hd__and2_1 _6294_ (.A(_2621_),
    .B(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__clkbuf_1 _6295_ (.A(_2623_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _6296_ (.A0(net10),
    .A1(_3403_),
    .S(_2596_),
    .X(_2624_));
 sky130_fd_sc_hd__and2_1 _6297_ (.A(_2624_),
    .B(_2622_),
    .X(_2625_));
 sky130_fd_sc_hd__clkbuf_1 _6298_ (.A(_2625_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _6299_ (.A0(net9),
    .A1(_3407_),
    .S(_2596_),
    .X(_2626_));
 sky130_fd_sc_hd__and2_1 _6300_ (.A(_2626_),
    .B(_2622_),
    .X(_2627_));
 sky130_fd_sc_hd__clkbuf_1 _6301_ (.A(_2627_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _6302_ (.A0(net8),
    .A1(_0693_),
    .S(_2596_),
    .X(_2628_));
 sky130_fd_sc_hd__and2_1 _6303_ (.A(_2628_),
    .B(_2622_),
    .X(_2629_));
 sky130_fd_sc_hd__clkbuf_1 _6304_ (.A(_2629_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _6305_ (.A0(net1),
    .A1(_0851_),
    .S(_2596_),
    .X(_2630_));
 sky130_fd_sc_hd__and2_1 _6306_ (.A(_2630_),
    .B(_2622_),
    .X(_2631_));
 sky130_fd_sc_hd__clkbuf_1 _6307_ (.A(_2631_),
    .X(_0184_));
 sky130_fd_sc_hd__or2_1 _6308_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .X(_2632_));
 sky130_fd_sc_hd__nand2_2 _6309_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2633_));
 sky130_fd_sc_hd__nand2_2 _6310_ (.A(_2632_),
    .B(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__o21ai_4 _6311_ (.A1(_3006_),
    .A2(_2634_),
    .B1(_2633_),
    .Y(_2635_));
 sky130_fd_sc_hd__or2_1 _6312_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .X(_2636_));
 sky130_fd_sc_hd__nand2_1 _6313_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2637_));
 sky130_fd_sc_hd__a21bo_2 _6314_ (.A1(_2635_),
    .A2(_2636_),
    .B1_N(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__or2_1 _6315_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .X(_2639_));
 sky130_fd_sc_hd__nand2_1 _6316_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2640_));
 sky130_fd_sc_hd__a21bo_2 _6317_ (.A1(_2638_),
    .A2(_2639_),
    .B1_N(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__and3_2 _6318_ (.A(_2641_),
    .B(\egd_top.BitStream_buffer.pc_previous[4] ),
    .C(\egd_top.BitStream_buffer.pc_previous[5] ),
    .X(_2642_));
 sky130_fd_sc_hd__xor2_4 _6319_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_2642_),
    .X(\egd_top.BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(_3036_),
    .B(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2643_));
 sky130_fd_sc_hd__inv_2 _6321_ (.A(_2643_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21oi_1 _6322_ (.A1(_2641_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[5] ),
    .Y(_2644_));
 sky130_fd_sc_hd__nor2_2 _6323_ (.A(_2644_),
    .B(_2642_),
    .Y(\egd_top.BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__nand2_1 _6324_ (.A(_3036_),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_2645_));
 sky130_fd_sc_hd__inv_2 _6325_ (.A(_2645_),
    .Y(_0182_));
 sky130_fd_sc_hd__xor2_4 _6326_ (.A(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B(_2641_),
    .X(\egd_top.BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__nand2_1 _6327_ (.A(_3036_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_2646_));
 sky130_fd_sc_hd__inv_2 _6328_ (.A(_2646_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_2 _6329_ (.A(_2639_),
    .B(_2640_),
    .Y(_2647_));
 sky130_fd_sc_hd__xnor2_4 _6330_ (.A(_2647_),
    .B(_2638_),
    .Y(\egd_top.BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__nand2_1 _6331_ (.A(_3036_),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2648_));
 sky130_fd_sc_hd__inv_2 _6332_ (.A(_2648_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_2 _6333_ (.A(_2636_),
    .B(_2637_),
    .Y(_2649_));
 sky130_fd_sc_hd__xnor2_4 _6334_ (.A(_2649_),
    .B(_2635_),
    .Y(\egd_top.BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__nand2_1 _6335_ (.A(_3036_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_2650_));
 sky130_fd_sc_hd__inv_2 _6336_ (.A(_2650_),
    .Y(_0179_));
 sky130_fd_sc_hd__xor2_4 _6337_ (.A(_3006_),
    .B(_2634_),
    .X(\egd_top.BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__nand2_1 _6338_ (.A(_3036_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2651_));
 sky130_fd_sc_hd__inv_2 _6339_ (.A(_2651_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_1 _6340_ (.A(_3008_),
    .B(_3036_),
    .Y(_2652_));
 sky130_fd_sc_hd__inv_2 _6341_ (.A(_2652_),
    .Y(_0177_));
 sky130_fd_sc_hd__or4b_1 _6342_ (.A(_3024_),
    .B(net198),
    .C(_3018_),
    .D_N(_3048_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_4 _6343_ (.A(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__clkbuf_4 _6344_ (.A(_2654_),
    .X(_2655_));
 sky130_fd_sc_hd__mux2_1 _6345_ (.A0(net7),
    .A1(_0637_),
    .S(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__and2_1 _6346_ (.A(_2656_),
    .B(_2622_),
    .X(_2657_));
 sky130_fd_sc_hd__clkbuf_1 _6347_ (.A(_2657_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _6348_ (.A0(net6),
    .A1(_0799_),
    .S(_2655_),
    .X(_2658_));
 sky130_fd_sc_hd__and2_1 _6349_ (.A(_2658_),
    .B(_2622_),
    .X(_2659_));
 sky130_fd_sc_hd__clkbuf_1 _6350_ (.A(_2659_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _6351_ (.A0(net5),
    .A1(_0661_),
    .S(_2655_),
    .X(_2660_));
 sky130_fd_sc_hd__and2_1 _6352_ (.A(_2660_),
    .B(_2622_),
    .X(_2661_));
 sky130_fd_sc_hd__clkbuf_1 _6353_ (.A(_2661_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _6354_ (.A0(net4),
    .A1(_3301_),
    .S(_2655_),
    .X(_2662_));
 sky130_fd_sc_hd__and2_1 _6355_ (.A(_2662_),
    .B(_2622_),
    .X(_2663_));
 sky130_fd_sc_hd__clkbuf_1 _6356_ (.A(_2663_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _6357_ (.A0(net3),
    .A1(_0663_),
    .S(_2655_),
    .X(_2664_));
 sky130_fd_sc_hd__and2_1 _6358_ (.A(_2664_),
    .B(_2622_),
    .X(_2665_));
 sky130_fd_sc_hd__clkbuf_1 _6359_ (.A(_2665_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _6360_ (.A0(net2),
    .A1(_0824_),
    .S(_2655_),
    .X(_2666_));
 sky130_fd_sc_hd__clkbuf_2 _6361_ (.A(net19),
    .X(_2667_));
 sky130_fd_sc_hd__and2_1 _6362_ (.A(_2666_),
    .B(_2667_),
    .X(_2668_));
 sky130_fd_sc_hd__clkbuf_1 _6363_ (.A(_2668_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _6364_ (.A0(net16),
    .A1(_0967_),
    .S(_2655_),
    .X(_2669_));
 sky130_fd_sc_hd__and2_1 _6365_ (.A(_2669_),
    .B(_2667_),
    .X(_2670_));
 sky130_fd_sc_hd__clkbuf_1 _6366_ (.A(_2670_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _6367_ (.A0(net15),
    .A1(_3323_),
    .S(_2655_),
    .X(_2671_));
 sky130_fd_sc_hd__and2_1 _6368_ (.A(_2671_),
    .B(_2667_),
    .X(_2672_));
 sky130_fd_sc_hd__clkbuf_1 _6369_ (.A(_2672_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _6370_ (.A0(net14),
    .A1(_0670_),
    .S(_2655_),
    .X(_2673_));
 sky130_fd_sc_hd__and2_1 _6371_ (.A(_2673_),
    .B(_2667_),
    .X(_2674_));
 sky130_fd_sc_hd__clkbuf_1 _6372_ (.A(_2674_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _6373_ (.A0(net13),
    .A1(_0831_),
    .S(_2655_),
    .X(_2675_));
 sky130_fd_sc_hd__and2_1 _6374_ (.A(_2675_),
    .B(_2667_),
    .X(_2676_));
 sky130_fd_sc_hd__clkbuf_1 _6375_ (.A(_2676_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _6376_ (.A0(net12),
    .A1(_3275_),
    .S(_2654_),
    .X(_2677_));
 sky130_fd_sc_hd__and2_1 _6377_ (.A(_2677_),
    .B(_2667_),
    .X(_2678_));
 sky130_fd_sc_hd__clkbuf_1 _6378_ (.A(_2678_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _6379_ (.A0(net11),
    .A1(_3282_),
    .S(_2654_),
    .X(_2679_));
 sky130_fd_sc_hd__and2_1 _6380_ (.A(_2679_),
    .B(_2667_),
    .X(_2680_));
 sky130_fd_sc_hd__clkbuf_1 _6381_ (.A(_2680_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _6382_ (.A0(net10),
    .A1(_0657_),
    .S(_2654_),
    .X(_2681_));
 sky130_fd_sc_hd__and2_1 _6383_ (.A(_2681_),
    .B(_2667_),
    .X(_2682_));
 sky130_fd_sc_hd__clkbuf_1 _6384_ (.A(_2682_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(net9),
    .A1(_0819_),
    .S(_2654_),
    .X(_2683_));
 sky130_fd_sc_hd__and2_1 _6386_ (.A(_2683_),
    .B(_2667_),
    .X(_2684_));
 sky130_fd_sc_hd__clkbuf_1 _6387_ (.A(_2684_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _6388_ (.A0(net8),
    .A1(_3326_),
    .S(_2654_),
    .X(_2685_));
 sky130_fd_sc_hd__and2_1 _6389_ (.A(_2685_),
    .B(_2667_),
    .X(_2686_));
 sky130_fd_sc_hd__clkbuf_1 _6390_ (.A(_2686_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _6391_ (.A0(net1),
    .A1(_3330_),
    .S(_2654_),
    .X(_2687_));
 sky130_fd_sc_hd__and2_1 _6392_ (.A(_2687_),
    .B(_3035_),
    .X(_2688_));
 sky130_fd_sc_hd__clkbuf_1 _6393_ (.A(_2688_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _6394_ (.A(net18),
    .B(net17),
    .Y(_2689_));
 sky130_fd_sc_hd__inv_2 _6395_ (.A(_2689_),
    .Y(_2690_));
 sky130_fd_sc_hd__and3b_1 _6396_ (.A_N(net21),
    .B(_2690_),
    .C(net20),
    .X(_2691_));
 sky130_fd_sc_hd__inv_2 _6397_ (.A(\egd_top.exp_golomb_decoding.te_range[2] ),
    .Y(_2692_));
 sky130_fd_sc_hd__and2_2 _6398_ (.A(_2691_),
    .B(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__nor2_1 _6399_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2694_));
 sky130_fd_sc_hd__nand2_1 _6400_ (.A(_2694_),
    .B(_3043_),
    .Y(_2695_));
 sky130_fd_sc_hd__nand2_1 _6401_ (.A(_1065_),
    .B(_1193_),
    .Y(_2696_));
 sky130_fd_sc_hd__nor2_1 _6402_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(_2696_),
    .Y(_2697_));
 sky130_fd_sc_hd__nand2_1 _6403_ (.A(_2697_),
    .B(_1318_),
    .Y(_2698_));
 sky130_fd_sc_hd__inv_2 _6404_ (.A(_2698_),
    .Y(_2699_));
 sky130_fd_sc_hd__and3_1 _6405_ (.A(_2699_),
    .B(_1442_),
    .C(_1566_),
    .X(_2700_));
 sky130_fd_sc_hd__inv_2 _6406_ (.A(_2700_),
    .Y(_2701_));
 sky130_fd_sc_hd__nor2_1 _6407_ (.A(_2695_),
    .B(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__nor2_1 _6408_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2703_));
 sky130_fd_sc_hd__inv_2 _6409_ (.A(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__nor2_1 _6410_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2704_),
    .Y(_2705_));
 sky130_fd_sc_hd__nand2_1 _6411_ (.A(_2705_),
    .B(_2049_),
    .Y(_2706_));
 sky130_fd_sc_hd__inv_2 _6412_ (.A(_2695_),
    .Y(_2707_));
 sky130_fd_sc_hd__nor2_1 _6413_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2708_));
 sky130_fd_sc_hd__nand2_2 _6414_ (.A(_2707_),
    .B(_2708_),
    .Y(_2709_));
 sky130_fd_sc_hd__a21o_1 _6415_ (.A1(_2700_),
    .A2(_2706_),
    .B1(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__nor2_2 _6416_ (.A(_2702_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__inv_6 _6417_ (.A(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__nand2_1 _6418_ (.A(_2287_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2713_));
 sky130_fd_sc_hd__nand2_1 _6419_ (.A(_2713_),
    .B(_2168_),
    .Y(_2714_));
 sky130_fd_sc_hd__nand2_1 _6420_ (.A(_2714_),
    .B(_2049_),
    .Y(_2715_));
 sky130_fd_sc_hd__nand2_1 _6421_ (.A(_2715_),
    .B(_1930_),
    .Y(_2716_));
 sky130_fd_sc_hd__nand2_1 _6422_ (.A(_2716_),
    .B(_1810_),
    .Y(_2717_));
 sky130_fd_sc_hd__nand2_1 _6423_ (.A(_2717_),
    .B(_1688_),
    .Y(_2718_));
 sky130_fd_sc_hd__nand2_1 _6424_ (.A(_2718_),
    .B(_1566_),
    .Y(_2719_));
 sky130_fd_sc_hd__nand2_1 _6425_ (.A(_2719_),
    .B(_1442_),
    .Y(_2720_));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(_2720_),
    .B(_2699_),
    .Y(_2721_));
 sky130_fd_sc_hd__a21oi_1 _6427_ (.A1(_1065_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2722_));
 sky130_fd_sc_hd__nand2_1 _6428_ (.A(_2721_),
    .B(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__nand2_2 _6429_ (.A(_2723_),
    .B(_2694_),
    .Y(_2724_));
 sky130_fd_sc_hd__o21ai_1 _6430_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_2049_),
    .Y(_2725_));
 sky130_fd_sc_hd__o211a_1 _6431_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .A2(_2725_),
    .B1(_1688_),
    .C1(_1810_),
    .X(_2726_));
 sky130_fd_sc_hd__a21o_1 _6432_ (.A1(_2698_),
    .A2(_2708_),
    .B1(_2695_),
    .X(_2727_));
 sky130_fd_sc_hd__o21bai_4 _6433_ (.A1(_2726_),
    .A2(_2701_),
    .B1_N(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__nor2_2 _6434_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_2729_));
 sky130_fd_sc_hd__nand3_1 _6435_ (.A(_2724_),
    .B(_2728_),
    .C(_2729_),
    .Y(_2730_));
 sky130_fd_sc_hd__nor2_1 _6436_ (.A(_2712_),
    .B(_2730_),
    .Y(_2731_));
 sky130_fd_sc_hd__inv_2 _6437_ (.A(_2731_),
    .Y(_2732_));
 sky130_fd_sc_hd__nor2_1 _6438_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .B(_2732_),
    .Y(_2733_));
 sky130_fd_sc_hd__inv_2 _6439_ (.A(_2728_),
    .Y(_2734_));
 sky130_fd_sc_hd__nor2_1 _6440_ (.A(_2734_),
    .B(_2712_),
    .Y(_2735_));
 sky130_fd_sc_hd__nand2_2 _6441_ (.A(_2724_),
    .B(_2729_),
    .Y(_2736_));
 sky130_fd_sc_hd__nand2_1 _6442_ (.A(_2735_),
    .B(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand2_1 _6443_ (.A(_2734_),
    .B(_2709_),
    .Y(_2738_));
 sky130_fd_sc_hd__inv_2 _6444_ (.A(_2738_),
    .Y(_2739_));
 sky130_fd_sc_hd__nand3_1 _6445_ (.A(_2739_),
    .B(_2736_),
    .C(_1193_),
    .Y(_2740_));
 sky130_fd_sc_hd__o21ai_1 _6446_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .A2(_2737_),
    .B1(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__nor2_1 _6447_ (.A(_2733_),
    .B(_2741_),
    .Y(_2742_));
 sky130_fd_sc_hd__nand3_4 _6448_ (.A(_2724_),
    .B(_2734_),
    .C(_2729_),
    .Y(_2743_));
 sky130_fd_sc_hd__inv_2 _6449_ (.A(_2743_),
    .Y(_2744_));
 sky130_fd_sc_hd__and3_1 _6450_ (.A(_2744_),
    .B(_1442_),
    .C(_2709_),
    .X(_2745_));
 sky130_fd_sc_hd__inv_2 _6451_ (.A(_2730_),
    .Y(_2746_));
 sky130_fd_sc_hd__and3_1 _6452_ (.A(_2746_),
    .B(_0931_),
    .C(_2709_),
    .X(_2747_));
 sky130_fd_sc_hd__nor2_1 _6453_ (.A(_2745_),
    .B(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__o21ai_1 _6454_ (.A1(_2712_),
    .A2(_2743_),
    .B1(_2168_),
    .Y(_2749_));
 sky130_fd_sc_hd__nor2_1 _6455_ (.A(_2712_),
    .B(_2743_),
    .Y(_2750_));
 sky130_fd_sc_hd__nand2_1 _6456_ (.A(_2750_),
    .B(_2406_),
    .Y(_2751_));
 sky130_fd_sc_hd__nand2_2 _6457_ (.A(_2749_),
    .B(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__nor2_2 _6458_ (.A(_2728_),
    .B(_2712_),
    .Y(_2753_));
 sky130_fd_sc_hd__nand2_1 _6459_ (.A(_2752_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__nand3_2 _6460_ (.A(_2742_),
    .B(_2748_),
    .C(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__clkbuf_4 _6461_ (.A(_3004_),
    .X(_2756_));
 sky130_fd_sc_hd__nand2_2 _6462_ (.A(_2755_),
    .B(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__inv_2 _6463_ (.A(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__or2_1 _6464_ (.A(_2693_),
    .B(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__inv_2 _6465_ (.A(_3004_),
    .Y(_2760_));
 sky130_fd_sc_hd__a311o_1 _6466_ (.A1(_2736_),
    .A2(_2710_),
    .A3(_2728_),
    .B1(_2760_),
    .C1(_2702_),
    .X(_2761_));
 sky130_fd_sc_hd__nand2_1 _6467_ (.A(_2761_),
    .B(_2693_),
    .Y(_2762_));
 sky130_fd_sc_hd__nor2_1 _6468_ (.A(net18),
    .B(_3003_),
    .Y(_2763_));
 sky130_fd_sc_hd__nand2_1 _6469_ (.A(_2744_),
    .B(_2711_),
    .Y(_2764_));
 sky130_fd_sc_hd__nand2_1 _6470_ (.A(_2764_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2765_));
 sky130_fd_sc_hd__buf_6 _6471_ (.A(_2750_),
    .X(_2766_));
 sky130_fd_sc_hd__nand2_1 _6472_ (.A(_2766_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2767_));
 sky130_fd_sc_hd__nand2_1 _6473_ (.A(_2765_),
    .B(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__o21ai_1 _6474_ (.A1(_2712_),
    .A2(_2743_),
    .B1(_2049_),
    .Y(_2769_));
 sky130_fd_sc_hd__nand3_1 _6475_ (.A(_2744_),
    .B(_2287_),
    .C(_2711_),
    .Y(_2770_));
 sky130_fd_sc_hd__nand2_1 _6476_ (.A(_2769_),
    .B(_2770_),
    .Y(_2771_));
 sky130_fd_sc_hd__nand2_1 _6477_ (.A(_2768_),
    .B(_2771_),
    .Y(_2772_));
 sky130_fd_sc_hd__o21ai_1 _6478_ (.A1(_2712_),
    .A2(_2743_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2773_));
 sky130_fd_sc_hd__nand3_1 _6479_ (.A(_2744_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .C(_2711_),
    .Y(_2774_));
 sky130_fd_sc_hd__nand2_1 _6480_ (.A(_2773_),
    .B(_2774_),
    .Y(_2775_));
 sky130_fd_sc_hd__nand2_1 _6481_ (.A(_2752_),
    .B(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__nand3_1 _6482_ (.A(_2772_),
    .B(_2776_),
    .C(_2753_),
    .Y(_2777_));
 sky130_fd_sc_hd__and2_1 _6483_ (.A(_2744_),
    .B(_2709_),
    .X(_2778_));
 sky130_fd_sc_hd__nor2_1 _6484_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2779_));
 sky130_fd_sc_hd__inv_2 _6485_ (.A(_2779_),
    .Y(_2780_));
 sky130_fd_sc_hd__nand2_1 _6486_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2781_));
 sky130_fd_sc_hd__nand2_1 _6487_ (.A(_2780_),
    .B(_2781_),
    .Y(_2782_));
 sky130_fd_sc_hd__nand2_1 _6488_ (.A(_2778_),
    .B(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__xnor2_1 _6489_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2784_));
 sky130_fd_sc_hd__nand3_1 _6490_ (.A(_2746_),
    .B(_2709_),
    .C(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(_2783_),
    .B(_2785_),
    .Y(_2786_));
 sky130_fd_sc_hd__xor2_1 _6492_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .X(_2787_));
 sky130_fd_sc_hd__nand2_1 _6493_ (.A(_2739_),
    .B(_2736_),
    .Y(_2788_));
 sky130_fd_sc_hd__nor2_2 _6494_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2789_));
 sky130_fd_sc_hd__inv_2 _6495_ (.A(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__nand2_1 _6496_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2791_));
 sky130_fd_sc_hd__nand2_1 _6497_ (.A(_2790_),
    .B(_2791_),
    .Y(_2792_));
 sky130_fd_sc_hd__nand3_1 _6498_ (.A(_2735_),
    .B(_2736_),
    .C(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__nand2_1 _6499_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2794_));
 sky130_fd_sc_hd__nand2_1 _6500_ (.A(_2704_),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__nand2_1 _6501_ (.A(_2731_),
    .B(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__o211ai_1 _6502_ (.A1(_2787_),
    .A2(_2788_),
    .B1(_2793_),
    .C1(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__nor2_1 _6503_ (.A(_2786_),
    .B(_2797_),
    .Y(_2798_));
 sky130_fd_sc_hd__nand2_1 _6504_ (.A(_2777_),
    .B(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__nand3_1 _6505_ (.A(_2799_),
    .B(_2756_),
    .C(_2755_),
    .Y(_2800_));
 sky130_fd_sc_hd__nor2_2 _6506_ (.A(net17),
    .B(_3002_),
    .Y(_2801_));
 sky130_fd_sc_hd__a22o_1 _6507_ (.A1(_2758_),
    .A2(_2763_),
    .B1(_2800_),
    .B2(_2801_),
    .X(_2802_));
 sky130_fd_sc_hd__nand2_2 _6508_ (.A(_2799_),
    .B(_2756_),
    .Y(_2803_));
 sky130_fd_sc_hd__nand2_1 _6509_ (.A(_2803_),
    .B(_2757_),
    .Y(_2804_));
 sky130_fd_sc_hd__a32o_2 _6510_ (.A1(_2690_),
    .A2(_2759_),
    .A3(_2762_),
    .B1(_2802_),
    .B2(_2804_),
    .X(net20));
 sky130_fd_sc_hd__a31o_1 _6511_ (.A1(_2691_),
    .A2(net18),
    .A3(_2692_),
    .B1(_3003_),
    .X(_2805_));
 sky130_fd_sc_hd__nand2_1 _6512_ (.A(_2752_),
    .B(_2771_),
    .Y(_2806_));
 sky130_fd_sc_hd__o21ai_1 _6513_ (.A1(_2712_),
    .A2(_2743_),
    .B1(_1930_),
    .Y(_2807_));
 sky130_fd_sc_hd__nand2_1 _6514_ (.A(_2750_),
    .B(_2168_),
    .Y(_2808_));
 sky130_fd_sc_hd__nand2_1 _6515_ (.A(_2807_),
    .B(_2808_),
    .Y(_2809_));
 sky130_fd_sc_hd__nand2_1 _6516_ (.A(_2806_),
    .B(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__o21ai_1 _6517_ (.A1(_2712_),
    .A2(_2743_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2811_));
 sky130_fd_sc_hd__nand2_1 _6518_ (.A(_2766_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2812_));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(_2811_),
    .B(_2812_),
    .Y(_2813_));
 sky130_fd_sc_hd__nand3_1 _6520_ (.A(_2752_),
    .B(_2813_),
    .C(_2771_),
    .Y(_2814_));
 sky130_fd_sc_hd__nand3_1 _6521_ (.A(_2810_),
    .B(_2814_),
    .C(_2753_),
    .Y(_2815_));
 sky130_fd_sc_hd__nor2_1 _6522_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2780_),
    .Y(_2816_));
 sky130_fd_sc_hd__nor2_1 _6523_ (.A(_1193_),
    .B(_2779_),
    .Y(_2817_));
 sky130_fd_sc_hd__o21ai_1 _6524_ (.A1(_2816_),
    .A2(_2817_),
    .B1(_2778_),
    .Y(_2818_));
 sky130_fd_sc_hd__nor2_1 _6525_ (.A(_1688_),
    .B(_2703_),
    .Y(_2819_));
 sky130_fd_sc_hd__o21ai_1 _6526_ (.A1(_2705_),
    .A2(_2819_),
    .B1(_2731_),
    .Y(_2820_));
 sky130_fd_sc_hd__nand2_1 _6527_ (.A(_2818_),
    .B(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__and2_1 _6528_ (.A(_2696_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .X(_2822_));
 sky130_fd_sc_hd__nor2_1 _6529_ (.A(_2697_),
    .B(_2822_),
    .Y(_2823_));
 sky130_fd_sc_hd__nor2_1 _6530_ (.A(_1442_),
    .B(_2789_),
    .Y(_2824_));
 sky130_fd_sc_hd__nor2_1 _6531_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2790_),
    .Y(_2825_));
 sky130_fd_sc_hd__inv_2 _6532_ (.A(_2737_),
    .Y(_2826_));
 sky130_fd_sc_hd__o21ai_1 _6533_ (.A1(_2824_),
    .A2(_2825_),
    .B1(_2826_),
    .Y(_2827_));
 sky130_fd_sc_hd__o21ai_1 _6534_ (.A1(_2788_),
    .A2(_2823_),
    .B1(_2827_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor2_1 _6535_ (.A(_2821_),
    .B(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__nand2_1 _6536_ (.A(_2815_),
    .B(_2829_),
    .Y(_2830_));
 sky130_fd_sc_hd__nand2_2 _6537_ (.A(_2830_),
    .B(_2756_),
    .Y(_2831_));
 sky130_fd_sc_hd__or2_1 _6538_ (.A(_2803_),
    .B(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__nand2_2 _6539_ (.A(_2831_),
    .B(_2803_),
    .Y(_2833_));
 sky130_fd_sc_hd__nand3_1 _6540_ (.A(_2832_),
    .B(_2833_),
    .C(_2801_),
    .Y(_2834_));
 sky130_fd_sc_hd__o21ai_4 _6541_ (.A1(_2803_),
    .A2(_2805_),
    .B1(_2834_),
    .Y(net21));
 sky130_fd_sc_hd__o21ai_1 _6542_ (.A1(_2803_),
    .A2(_2831_),
    .B1(_2758_),
    .Y(_2835_));
 sky130_fd_sc_hd__nand2_1 _6543_ (.A(_2835_),
    .B(_2833_),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_1 _6544_ (.A(_2775_),
    .B(_2768_),
    .Y(_2837_));
 sky130_fd_sc_hd__nand2_1 _6545_ (.A(_2766_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2838_));
 sky130_fd_sc_hd__o21ai_1 _6546_ (.A1(_1810_),
    .A2(_2766_),
    .B1(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__nand3_1 _6547_ (.A(_2837_),
    .B(_2839_),
    .C(_2809_),
    .Y(_2840_));
 sky130_fd_sc_hd__nand3_1 _6548_ (.A(_2752_),
    .B(_2809_),
    .C(_2771_),
    .Y(_2841_));
 sky130_fd_sc_hd__nand2_1 _6549_ (.A(_2766_),
    .B(_2049_),
    .Y(_2842_));
 sky130_fd_sc_hd__o21ai_1 _6550_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .A2(_2766_),
    .B1(_2842_),
    .Y(_2843_));
 sky130_fd_sc_hd__nand2_1 _6551_ (.A(_2841_),
    .B(_2843_),
    .Y(_2844_));
 sky130_fd_sc_hd__nand3_1 _6552_ (.A(_2840_),
    .B(_2844_),
    .C(_2753_),
    .Y(_2845_));
 sky130_fd_sc_hd__nand2_1 _6553_ (.A(_2816_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2846_));
 sky130_fd_sc_hd__or2_1 _6554_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(_2816_),
    .X(_2847_));
 sky130_fd_sc_hd__and3_1 _6555_ (.A(_2778_),
    .B(_2846_),
    .C(_2847_),
    .X(_2848_));
 sky130_fd_sc_hd__or2_1 _6556_ (.A(_1566_),
    .B(_2705_),
    .X(_2849_));
 sky130_fd_sc_hd__nor2_1 _6557_ (.A(_2704_),
    .B(_2790_),
    .Y(_2850_));
 sky130_fd_sc_hd__inv_2 _6558_ (.A(_2850_),
    .Y(_2851_));
 sky130_fd_sc_hd__nand2_1 _6559_ (.A(_2849_),
    .B(_2851_),
    .Y(_2852_));
 sky130_fd_sc_hd__mux2_1 _6560_ (.A0(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .A1(_2782_),
    .S(_2789_),
    .X(_2853_));
 sky130_fd_sc_hd__a22o_1 _6561_ (.A1(_2731_),
    .A2(_2852_),
    .B1(_2826_),
    .B2(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__nor2_1 _6562_ (.A(_2848_),
    .B(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__a21oi_1 _6563_ (.A1(_2845_),
    .A2(_2855_),
    .B1(_2760_),
    .Y(_2856_));
 sky130_fd_sc_hd__nand2_1 _6564_ (.A(_2836_),
    .B(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__nand2_1 _6565_ (.A(_2845_),
    .B(_2855_),
    .Y(_2858_));
 sky130_fd_sc_hd__nand2_1 _6566_ (.A(_2858_),
    .B(_2756_),
    .Y(_2859_));
 sky130_fd_sc_hd__nand3_1 _6567_ (.A(_2835_),
    .B(_2833_),
    .C(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__nand2_1 _6568_ (.A(_2857_),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__nand2_1 _6569_ (.A(_2861_),
    .B(_2801_),
    .Y(_2862_));
 sky130_fd_sc_hd__or2_1 _6570_ (.A(_2805_),
    .B(_2831_),
    .X(_2863_));
 sky130_fd_sc_hd__nand2_1 _6571_ (.A(net20),
    .B(net21),
    .Y(_2864_));
 sky130_fd_sc_hd__a21oi_1 _6572_ (.A1(_2862_),
    .A2(_2863_),
    .B1(_2864_),
    .Y(_2865_));
 sky130_fd_sc_hd__nand3_1 _6573_ (.A(_2862_),
    .B(_2864_),
    .C(_2863_),
    .Y(_2866_));
 sky130_fd_sc_hd__nand2_1 _6574_ (.A(_2866_),
    .B(_2690_),
    .Y(_2867_));
 sky130_fd_sc_hd__nor2_1 _6575_ (.A(_2865_),
    .B(_2867_),
    .Y(\egd_top.exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__or3_1 _6576_ (.A(_2760_),
    .B(_2693_),
    .C(_2736_),
    .X(_2868_));
 sky130_fd_sc_hd__inv_2 _6577_ (.A(_2868_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__or3_1 _6578_ (.A(_2760_),
    .B(_2693_),
    .C(_2728_),
    .X(_2869_));
 sky130_fd_sc_hd__inv_2 _6579_ (.A(_2869_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__or3_1 _6580_ (.A(_2760_),
    .B(_2693_),
    .C(_2710_),
    .X(_2870_));
 sky130_fd_sc_hd__inv_2 _6581_ (.A(_2870_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__nand2_1 _6582_ (.A(_2862_),
    .B(_2863_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_1 _6583_ (.A(_2843_),
    .B(_2809_),
    .Y(_2871_));
 sky130_fd_sc_hd__nand2_1 _6584_ (.A(_2766_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2872_));
 sky130_fd_sc_hd__o21ai_2 _6585_ (.A1(_1688_),
    .A2(_2766_),
    .B1(_2872_),
    .Y(_2873_));
 sky130_fd_sc_hd__inv_2 _6586_ (.A(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__o21ai_1 _6587_ (.A1(_2806_),
    .A2(_2871_),
    .B1(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__nor2_1 _6588_ (.A(_2806_),
    .B(_2871_),
    .Y(_2876_));
 sky130_fd_sc_hd__nand2_1 _6589_ (.A(_2876_),
    .B(_2873_),
    .Y(_2877_));
 sky130_fd_sc_hd__nand3_1 _6590_ (.A(_2875_),
    .B(_2877_),
    .C(_2753_),
    .Y(_2878_));
 sky130_fd_sc_hd__nor2_1 _6591_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2850_),
    .Y(_2879_));
 sky130_fd_sc_hd__nor2_1 _6592_ (.A(_1442_),
    .B(_2851_),
    .Y(_2880_));
 sky130_fd_sc_hd__nand2_1 _6593_ (.A(_2789_),
    .B(_2779_),
    .Y(_2881_));
 sky130_fd_sc_hd__xor2_1 _6594_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__o32a_1 _6595_ (.A1(_2879_),
    .A2(_2880_),
    .A3(_2732_),
    .B1(_2737_),
    .B2(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__nand2_1 _6596_ (.A(_2878_),
    .B(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__nand2_2 _6597_ (.A(_2884_),
    .B(_2756_),
    .Y(_2885_));
 sky130_fd_sc_hd__nor2_1 _6598_ (.A(_2833_),
    .B(_2856_),
    .Y(_2886_));
 sky130_fd_sc_hd__nor2_1 _6599_ (.A(_2885_),
    .B(_2886_),
    .Y(_2887_));
 sky130_fd_sc_hd__nand2_1 _6600_ (.A(_2885_),
    .B(_2859_),
    .Y(_2888_));
 sky130_fd_sc_hd__nor2_1 _6601_ (.A(_2833_),
    .B(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__o21a_1 _6602_ (.A1(_2887_),
    .A2(_2889_),
    .B1(_2757_),
    .X(_2890_));
 sky130_fd_sc_hd__nor2_1 _6603_ (.A(_2800_),
    .B(_2831_),
    .Y(_2891_));
 sky130_fd_sc_hd__nand2_1 _6604_ (.A(_2856_),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__nor2_1 _6605_ (.A(_2885_),
    .B(_2892_),
    .Y(_2893_));
 sky130_fd_sc_hd__and2_1 _6606_ (.A(_2892_),
    .B(_2885_),
    .X(_2894_));
 sky130_fd_sc_hd__o21ai_1 _6607_ (.A1(_2893_),
    .A2(_2894_),
    .B1(_2758_),
    .Y(_2895_));
 sky130_fd_sc_hd__nand2_1 _6608_ (.A(_2895_),
    .B(_2801_),
    .Y(_2896_));
 sky130_fd_sc_hd__inv_2 _6609_ (.A(_2805_),
    .Y(_2897_));
 sky130_fd_sc_hd__nand2_1 _6610_ (.A(_2858_),
    .B(_2897_),
    .Y(_2898_));
 sky130_fd_sc_hd__o21ai_2 _6611_ (.A1(_2890_),
    .A2(_2896_),
    .B1(_2898_),
    .Y(net23));
 sky130_fd_sc_hd__nand2_1 _6612_ (.A(_2889_),
    .B(_2757_),
    .Y(_2899_));
 sky130_fd_sc_hd__o21ai_1 _6613_ (.A1(_2885_),
    .A2(_2892_),
    .B1(_2758_),
    .Y(_2900_));
 sky130_fd_sc_hd__nand2_1 _6614_ (.A(_2899_),
    .B(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__nor2_1 _6615_ (.A(_2813_),
    .B(_2839_),
    .Y(_2902_));
 sky130_fd_sc_hd__nand3_1 _6616_ (.A(_2902_),
    .B(_2837_),
    .C(_2874_),
    .Y(_2903_));
 sky130_fd_sc_hd__a21oi_1 _6617_ (.A1(_2766_),
    .A2(_1810_),
    .B1(_1566_),
    .Y(_2904_));
 sky130_fd_sc_hd__inv_2 _6618_ (.A(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__nand2_1 _6619_ (.A(_2903_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__nand3_1 _6620_ (.A(_2876_),
    .B(_2904_),
    .C(_2874_),
    .Y(_2907_));
 sky130_fd_sc_hd__nand3_1 _6621_ (.A(_2906_),
    .B(_2907_),
    .C(_2753_),
    .Y(_2908_));
 sky130_fd_sc_hd__nor2_1 _6622_ (.A(_2782_),
    .B(_2851_),
    .Y(_2909_));
 sky130_fd_sc_hd__a211o_1 _6623_ (.A1(_1318_),
    .A2(_2851_),
    .B1(_2909_),
    .C1(_2732_),
    .X(_2910_));
 sky130_fd_sc_hd__nand2_1 _6624_ (.A(_2908_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__nand2_1 _6625_ (.A(_2911_),
    .B(_2756_),
    .Y(_2912_));
 sky130_fd_sc_hd__nand2_1 _6626_ (.A(_2901_),
    .B(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__inv_2 _6627_ (.A(_2912_),
    .Y(_2914_));
 sky130_fd_sc_hd__nand3_1 _6628_ (.A(_2899_),
    .B(_2900_),
    .C(_2914_),
    .Y(_2915_));
 sky130_fd_sc_hd__nand3_1 _6629_ (.A(_2913_),
    .B(_2915_),
    .C(_2801_),
    .Y(_2916_));
 sky130_fd_sc_hd__nand2_1 _6630_ (.A(_2884_),
    .B(_2897_),
    .Y(_2917_));
 sky130_fd_sc_hd__nand2_1 _6631_ (.A(_2916_),
    .B(_2917_),
    .Y(net24));
 sky130_fd_sc_hd__nand3_1 _6632_ (.A(_2911_),
    .B(_2756_),
    .C(_2884_),
    .Y(_2918_));
 sky130_fd_sc_hd__inv_2 _6633_ (.A(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__nor3_1 _6634_ (.A(_2831_),
    .B(_2800_),
    .C(_2859_),
    .Y(_2920_));
 sky130_fd_sc_hd__nand2_1 _6635_ (.A(_2919_),
    .B(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__nor2_1 _6636_ (.A(_2904_),
    .B(_2873_),
    .Y(_2922_));
 sky130_fd_sc_hd__nand2_1 _6637_ (.A(_2876_),
    .B(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__o21ai_2 _6638_ (.A1(_1688_),
    .A2(_2764_),
    .B1(_1442_),
    .Y(_2924_));
 sky130_fd_sc_hd__inv_2 _6639_ (.A(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__nand2_1 _6640_ (.A(_2923_),
    .B(_2925_),
    .Y(_2926_));
 sky130_fd_sc_hd__nand3_1 _6641_ (.A(_2876_),
    .B(_2922_),
    .C(_2924_),
    .Y(_2927_));
 sky130_fd_sc_hd__nand3_1 _6642_ (.A(_2926_),
    .B(_2753_),
    .C(_2927_),
    .Y(_2928_));
 sky130_fd_sc_hd__nor2_2 _6643_ (.A(_2760_),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__inv_2 _6644_ (.A(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(_2921_),
    .B(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__nand3_1 _6646_ (.A(_2919_),
    .B(_2920_),
    .C(_2929_),
    .Y(_2932_));
 sky130_fd_sc_hd__nand2_1 _6647_ (.A(_2931_),
    .B(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__nand2_1 _6648_ (.A(_2933_),
    .B(_2758_),
    .Y(_2934_));
 sky130_fd_sc_hd__nand3_1 _6649_ (.A(_2886_),
    .B(_2885_),
    .C(_2912_),
    .Y(_2935_));
 sky130_fd_sc_hd__nand2_1 _6650_ (.A(_2935_),
    .B(_2929_),
    .Y(_2936_));
 sky130_fd_sc_hd__a21oi_1 _6651_ (.A1(_2911_),
    .A2(_2756_),
    .B1(_2929_),
    .Y(_2937_));
 sky130_fd_sc_hd__nand2_1 _6652_ (.A(_2889_),
    .B(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__nand2_1 _6653_ (.A(_2936_),
    .B(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__nand2_1 _6654_ (.A(_2939_),
    .B(_2757_),
    .Y(_2940_));
 sky130_fd_sc_hd__nand3_1 _6655_ (.A(_2934_),
    .B(_2940_),
    .C(_2801_),
    .Y(_2941_));
 sky130_fd_sc_hd__nand2_1 _6656_ (.A(_2911_),
    .B(_2897_),
    .Y(_2942_));
 sky130_fd_sc_hd__nand2_1 _6657_ (.A(_2941_),
    .B(_2942_),
    .Y(net25));
 sky130_fd_sc_hd__nand3_1 _6658_ (.A(_2893_),
    .B(_2929_),
    .C(_2914_),
    .Y(_2943_));
 sky130_fd_sc_hd__or2_1 _6659_ (.A(_2924_),
    .B(_2923_),
    .X(_2944_));
 sky130_fd_sc_hd__nand2_1 _6660_ (.A(_2944_),
    .B(_2766_),
    .Y(_2945_));
 sky130_fd_sc_hd__inv_2 _6661_ (.A(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__nand2_1 _6662_ (.A(_2946_),
    .B(_2756_),
    .Y(_2947_));
 sky130_fd_sc_hd__nand2_1 _6663_ (.A(_2943_),
    .B(_2947_),
    .Y(_2948_));
 sky130_fd_sc_hd__nand2_1 _6664_ (.A(_2948_),
    .B(_2758_),
    .Y(_2949_));
 sky130_fd_sc_hd__inv_2 _6665_ (.A(_2947_),
    .Y(_2950_));
 sky130_fd_sc_hd__nand2_1 _6666_ (.A(_2938_),
    .B(_2950_),
    .Y(_2951_));
 sky130_fd_sc_hd__nor2_1 _6667_ (.A(_2761_),
    .B(_2755_),
    .Y(_2952_));
 sky130_fd_sc_hd__nand2_1 _6668_ (.A(_2951_),
    .B(_2952_),
    .Y(_2953_));
 sky130_fd_sc_hd__nand2_1 _6669_ (.A(_2949_),
    .B(_2953_),
    .Y(_2954_));
 sky130_fd_sc_hd__nand2_1 _6670_ (.A(_2954_),
    .B(_2801_),
    .Y(_2955_));
 sky130_fd_sc_hd__a211o_1 _6671_ (.A1(net18),
    .A2(_2693_),
    .B1(_3003_),
    .C1(_2928_),
    .X(_2956_));
 sky130_fd_sc_hd__nand2_1 _6672_ (.A(_2955_),
    .B(_2956_),
    .Y(net26));
 sky130_fd_sc_hd__a211o_1 _6673_ (.A1(net18),
    .A2(_2693_),
    .B1(_3003_),
    .C1(_2945_),
    .X(_2957_));
 sky130_fd_sc_hd__a21bo_1 _6674_ (.A1(_2801_),
    .A2(_2952_),
    .B1_N(_2957_),
    .X(net27));
 sky130_fd_sc_hd__buf_1 _6675_ (.A(wb_clk_i),
    .X(_2958_));
 sky130_fd_sc_hd__buf_1 _6676_ (.A(clknet_1_1__leaf__2958_),
    .X(_2959_));
 sky130_fd_sc_hd__buf_1 _6677_ (.A(clknet_1_0__leaf__2959_),
    .X(_2960_));
 sky130_fd_sc_hd__inv_2 _6678__72 (.A(clknet_1_0__leaf__2960_),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _6679__73 (.A(clknet_1_0__leaf__2960_),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _6680__74 (.A(clknet_1_0__leaf__2960_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _6681__75 (.A(clknet_1_0__leaf__2960_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _6682__76 (.A(clknet_1_1__leaf__2960_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _6683__77 (.A(clknet_1_1__leaf__2960_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _6684__78 (.A(clknet_1_1__leaf__2960_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _6685__79 (.A(clknet_1_1__leaf__2960_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _6686__80 (.A(clknet_1_1__leaf__2960_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _6687__81 (.A(clknet_1_1__leaf__2960_),
    .Y(net115));
 sky130_fd_sc_hd__buf_1 _6688_ (.A(clknet_1_0__leaf__2959_),
    .X(_2961_));
 sky130_fd_sc_hd__inv_2 _6689__82 (.A(clknet_1_1__leaf__2961_),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _6690__83 (.A(clknet_1_1__leaf__2961_),
    .Y(net117));
 sky130_fd_sc_hd__inv_2 _6691__84 (.A(clknet_1_1__leaf__2961_),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _6692__85 (.A(clknet_1_1__leaf__2961_),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _6693__86 (.A(clknet_1_1__leaf__2961_),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _6694__87 (.A(clknet_1_1__leaf__2961_),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _6695__88 (.A(clknet_1_0__leaf__2961_),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _6696__89 (.A(clknet_1_0__leaf__2961_),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _6697__90 (.A(clknet_1_0__leaf__2961_),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _6698__91 (.A(clknet_1_0__leaf__2961_),
    .Y(net125));
 sky130_fd_sc_hd__buf_1 _6699_ (.A(clknet_1_0__leaf__2959_),
    .X(_2962_));
 sky130_fd_sc_hd__inv_2 _6700__92 (.A(clknet_1_1__leaf__2962_),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _6701__93 (.A(clknet_1_1__leaf__2962_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _6702__94 (.A(clknet_1_1__leaf__2962_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _6703__95 (.A(clknet_1_1__leaf__2962_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _6704__96 (.A(clknet_1_0__leaf__2962_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _6705__97 (.A(clknet_1_0__leaf__2962_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _6706__98 (.A(clknet_1_0__leaf__2962_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _6707__99 (.A(clknet_1_0__leaf__2962_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _6708__100 (.A(clknet_1_0__leaf__2962_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _6709__101 (.A(clknet_1_0__leaf__2962_),
    .Y(net135));
 sky130_fd_sc_hd__buf_1 _6710_ (.A(clknet_1_0__leaf__2959_),
    .X(_2963_));
 sky130_fd_sc_hd__inv_2 _6711__102 (.A(clknet_1_1__leaf__2963_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _6712__103 (.A(clknet_1_0__leaf__2963_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _6713__104 (.A(clknet_1_0__leaf__2963_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _6714__105 (.A(clknet_1_0__leaf__2963_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _6715__106 (.A(clknet_1_0__leaf__2963_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _6716__107 (.A(clknet_1_1__leaf__2963_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _6717__108 (.A(clknet_1_1__leaf__2963_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _6718__109 (.A(clknet_1_1__leaf__2963_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _6719__110 (.A(clknet_1_1__leaf__2963_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _6720__111 (.A(clknet_1_1__leaf__2963_),
    .Y(net145));
 sky130_fd_sc_hd__buf_1 _6721_ (.A(clknet_1_1__leaf__2959_),
    .X(_2964_));
 sky130_fd_sc_hd__inv_2 _6722__112 (.A(clknet_1_0__leaf__2964_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _6723__113 (.A(clknet_1_0__leaf__2964_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _6724__114 (.A(clknet_1_0__leaf__2964_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _6725__115 (.A(clknet_1_0__leaf__2964_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _6726__116 (.A(clknet_1_0__leaf__2964_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _6727__117 (.A(clknet_1_1__leaf__2964_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _6728__118 (.A(clknet_1_1__leaf__2964_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _6729__119 (.A(clknet_1_1__leaf__2964_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _6730__120 (.A(clknet_1_1__leaf__2964_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _6731__121 (.A(clknet_1_1__leaf__2964_),
    .Y(net155));
 sky130_fd_sc_hd__buf_1 _6732_ (.A(clknet_1_1__leaf__2959_),
    .X(_2965_));
 sky130_fd_sc_hd__inv_2 _6733__122 (.A(clknet_1_0__leaf__2965_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _6734__123 (.A(clknet_1_0__leaf__2965_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _6735__124 (.A(clknet_1_0__leaf__2965_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _6736__125 (.A(clknet_1_0__leaf__2965_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _6737__126 (.A(clknet_1_0__leaf__2965_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _6738__127 (.A(clknet_1_0__leaf__2965_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _6739__128 (.A(clknet_1_1__leaf__2965_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _6740__129 (.A(clknet_1_1__leaf__2965_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _6741__130 (.A(clknet_1_1__leaf__2965_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _6742__131 (.A(clknet_1_1__leaf__2965_),
    .Y(net165));
 sky130_fd_sc_hd__buf_1 _6743_ (.A(clknet_1_1__leaf__2959_),
    .X(_2966_));
 sky130_fd_sc_hd__inv_2 _6744__132 (.A(clknet_1_0__leaf__2966_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _6745__133 (.A(clknet_1_0__leaf__2966_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _6746__134 (.A(clknet_1_0__leaf__2966_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _6747__135 (.A(clknet_1_0__leaf__2966_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _6748__136 (.A(clknet_1_0__leaf__2966_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _6749__137 (.A(clknet_1_1__leaf__2966_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _6750__138 (.A(clknet_1_1__leaf__2966_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _6751__139 (.A(clknet_1_1__leaf__2966_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _6752__140 (.A(clknet_1_1__leaf__2966_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _6753__141 (.A(clknet_1_1__leaf__2966_),
    .Y(net175));
 sky130_fd_sc_hd__buf_1 _6754_ (.A(clknet_1_1__leaf__2959_),
    .X(_2967_));
 sky130_fd_sc_hd__inv_2 _6755__142 (.A(clknet_1_1__leaf__2967_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _6756__143 (.A(clknet_1_1__leaf__2967_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _6757__144 (.A(clknet_1_1__leaf__2967_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _6758__145 (.A(clknet_1_1__leaf__2967_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _6759__146 (.A(clknet_1_1__leaf__2967_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _6760__147 (.A(clknet_1_0__leaf__2967_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _6761__148 (.A(clknet_1_0__leaf__2967_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _6762__149 (.A(clknet_1_0__leaf__2967_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _6763__150 (.A(clknet_1_0__leaf__2967_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _6764__151 (.A(clknet_1_0__leaf__2967_),
    .Y(net185));
 sky130_fd_sc_hd__buf_1 _6765_ (.A(clknet_1_1__leaf__2959_),
    .X(_2968_));
 sky130_fd_sc_hd__inv_2 _6766__152 (.A(clknet_1_1__leaf__2968_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _6767__153 (.A(clknet_1_1__leaf__2968_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _6768__154 (.A(clknet_1_1__leaf__2968_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _6769__155 (.A(clknet_1_1__leaf__2968_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _6770__156 (.A(clknet_1_0__leaf__2968_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _6771__157 (.A(clknet_1_1__leaf__2968_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _6772__158 (.A(clknet_1_0__leaf__2968_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _6773__159 (.A(clknet_1_0__leaf__2968_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _6774__160 (.A(clknet_1_0__leaf__2968_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _6775__161 (.A(clknet_1_0__leaf__2968_),
    .Y(net195));
 sky130_fd_sc_hd__buf_1 _6776_ (.A(clknet_1_1__leaf__2958_),
    .X(_2969_));
 sky130_fd_sc_hd__inv_2 _6777__2 (.A(clknet_1_1__leaf__2969_),
    .Y(net36));
 sky130_fd_sc_hd__inv_2 _6778__3 (.A(clknet_1_1__leaf__2969_),
    .Y(net37));
 sky130_fd_sc_hd__inv_2 _6779__4 (.A(clknet_1_1__leaf__2969_),
    .Y(net38));
 sky130_fd_sc_hd__inv_2 _6780__5 (.A(clknet_1_1__leaf__2969_),
    .Y(net39));
 sky130_fd_sc_hd__inv_2 _6781__6 (.A(clknet_1_0__leaf__2969_),
    .Y(net40));
 sky130_fd_sc_hd__inv_2 _6782__7 (.A(clknet_1_1__leaf__2969_),
    .Y(net41));
 sky130_fd_sc_hd__inv_2 _6783__8 (.A(clknet_1_0__leaf__2969_),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _6784__9 (.A(clknet_1_0__leaf__2969_),
    .Y(net43));
 sky130_fd_sc_hd__inv_2 _6785__10 (.A(clknet_1_0__leaf__2969_),
    .Y(net44));
 sky130_fd_sc_hd__inv_2 _6786__11 (.A(clknet_1_0__leaf__2969_),
    .Y(net45));
 sky130_fd_sc_hd__buf_1 _6787_ (.A(clknet_1_1__leaf__2958_),
    .X(_2970_));
 sky130_fd_sc_hd__inv_2 _6788__12 (.A(clknet_1_1__leaf__2970_),
    .Y(net46));
 sky130_fd_sc_hd__inv_2 _6789__13 (.A(clknet_1_1__leaf__2970_),
    .Y(net47));
 sky130_fd_sc_hd__inv_2 _6790__14 (.A(clknet_1_1__leaf__2970_),
    .Y(net48));
 sky130_fd_sc_hd__inv_2 _6791__15 (.A(clknet_1_1__leaf__2970_),
    .Y(net49));
 sky130_fd_sc_hd__inv_2 _6792__16 (.A(clknet_1_1__leaf__2970_),
    .Y(net50));
 sky130_fd_sc_hd__inv_2 _6793__17 (.A(clknet_1_0__leaf__2970_),
    .Y(net51));
 sky130_fd_sc_hd__inv_2 _6794__18 (.A(clknet_1_0__leaf__2970_),
    .Y(net52));
 sky130_fd_sc_hd__inv_2 _6795__19 (.A(clknet_1_0__leaf__2970_),
    .Y(net53));
 sky130_fd_sc_hd__inv_2 _6796__20 (.A(clknet_1_0__leaf__2970_),
    .Y(net54));
 sky130_fd_sc_hd__inv_2 _6797__21 (.A(clknet_1_0__leaf__2970_),
    .Y(net55));
 sky130_fd_sc_hd__buf_1 _6798_ (.A(clknet_1_0__leaf__2958_),
    .X(_2971_));
 sky130_fd_sc_hd__inv_2 _6799__22 (.A(clknet_1_1__leaf__2971_),
    .Y(net56));
 sky130_fd_sc_hd__inv_2 _6800__23 (.A(clknet_1_1__leaf__2971_),
    .Y(net57));
 sky130_fd_sc_hd__inv_2 _6801__24 (.A(clknet_1_1__leaf__2971_),
    .Y(net58));
 sky130_fd_sc_hd__inv_2 _6802__25 (.A(clknet_1_1__leaf__2971_),
    .Y(net59));
 sky130_fd_sc_hd__inv_2 _6803__26 (.A(clknet_1_1__leaf__2971_),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 _6804__27 (.A(clknet_1_0__leaf__2971_),
    .Y(net61));
 sky130_fd_sc_hd__inv_2 _6805__28 (.A(clknet_1_0__leaf__2971_),
    .Y(net62));
 sky130_fd_sc_hd__inv_2 _6806__29 (.A(clknet_1_0__leaf__2971_),
    .Y(net63));
 sky130_fd_sc_hd__inv_2 _6807__30 (.A(clknet_1_0__leaf__2971_),
    .Y(net64));
 sky130_fd_sc_hd__inv_2 _6808__31 (.A(clknet_1_0__leaf__2971_),
    .Y(net65));
 sky130_fd_sc_hd__buf_1 _6809_ (.A(clknet_1_0__leaf__2958_),
    .X(_2972_));
 sky130_fd_sc_hd__inv_2 _6810__32 (.A(clknet_1_0__leaf__2972_),
    .Y(net66));
 sky130_fd_sc_hd__inv_2 _6811__33 (.A(clknet_1_0__leaf__2972_),
    .Y(net67));
 sky130_fd_sc_hd__inv_2 _6812__34 (.A(clknet_1_0__leaf__2972_),
    .Y(net68));
 sky130_fd_sc_hd__inv_2 _6813__35 (.A(clknet_1_0__leaf__2972_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _6814__36 (.A(clknet_1_0__leaf__2972_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _6815__37 (.A(clknet_1_0__leaf__2972_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _6816__38 (.A(clknet_1_1__leaf__2972_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _6817__39 (.A(clknet_1_1__leaf__2972_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _6818__40 (.A(clknet_1_1__leaf__2972_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _6819__41 (.A(clknet_1_1__leaf__2972_),
    .Y(net75));
 sky130_fd_sc_hd__buf_1 _6820_ (.A(clknet_1_1__leaf__2958_),
    .X(_2973_));
 sky130_fd_sc_hd__inv_2 _6821__42 (.A(clknet_1_0__leaf__2973_),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _6822__43 (.A(clknet_1_0__leaf__2973_),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _6823__44 (.A(clknet_1_0__leaf__2973_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _6824__45 (.A(clknet_1_0__leaf__2973_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _6825__46 (.A(clknet_1_0__leaf__2973_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _6826__47 (.A(clknet_1_1__leaf__2973_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _6827__48 (.A(clknet_1_0__leaf__2973_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _6828__49 (.A(clknet_1_1__leaf__2973_),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _6829__50 (.A(clknet_1_1__leaf__2973_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _6830__51 (.A(clknet_1_1__leaf__2973_),
    .Y(net85));
 sky130_fd_sc_hd__buf_1 _6831_ (.A(clknet_1_0__leaf__2958_),
    .X(_2974_));
 sky130_fd_sc_hd__inv_2 _6832__52 (.A(clknet_1_1__leaf__2974_),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _6833__53 (.A(clknet_1_1__leaf__2974_),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _6834__54 (.A(clknet_1_1__leaf__2974_),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _6835__55 (.A(clknet_1_1__leaf__2974_),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _6836__56 (.A(clknet_1_1__leaf__2974_),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _6837__57 (.A(clknet_1_0__leaf__2974_),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _6838__58 (.A(clknet_1_0__leaf__2974_),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _6839__59 (.A(clknet_1_0__leaf__2974_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _6840__60 (.A(clknet_1_0__leaf__2974_),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _6841__61 (.A(clknet_1_0__leaf__2974_),
    .Y(net95));
 sky130_fd_sc_hd__buf_1 _6842_ (.A(clknet_1_0__leaf__2958_),
    .X(_2975_));
 sky130_fd_sc_hd__inv_2 _6843__62 (.A(clknet_1_1__leaf__2975_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _6844__63 (.A(clknet_1_1__leaf__2975_),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _6845__64 (.A(clknet_1_1__leaf__2975_),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _6846__65 (.A(clknet_1_1__leaf__2975_),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _6847__66 (.A(clknet_1_0__leaf__2975_),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _6848__67 (.A(clknet_1_0__leaf__2975_),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _6849__68 (.A(clknet_1_0__leaf__2975_),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _6850__69 (.A(clknet_1_0__leaf__2975_),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _6851__70 (.A(clknet_1_0__leaf__2975_),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _6852__71 (.A(clknet_1_0__leaf__2975_),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _6853__1 (.A(clknet_1_0__leaf__2959_),
    .Y(net35));
 sky130_fd_sc_hd__dfxtp_1 _6854_ (.CLK(net106),
    .D(_0161_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfxtp_1 _6855_ (.CLK(net107),
    .D(_0162_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfxtp_1 _6856_ (.CLK(net108),
    .D(_0163_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfxtp_1 _6857_ (.CLK(net109),
    .D(_0164_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfxtp_1 _6858_ (.CLK(net110),
    .D(_0165_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfxtp_1 _6859_ (.CLK(net111),
    .D(_0166_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfxtp_1 _6860_ (.CLK(net112),
    .D(_0167_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfxtp_1 _6861_ (.CLK(net113),
    .D(_0168_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfxtp_1 _6862_ (.CLK(net114),
    .D(_0169_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfxtp_1 _6863_ (.CLK(net115),
    .D(_0170_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfxtp_1 _6864_ (.CLK(net116),
    .D(_0171_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfxtp_1 _6865_ (.CLK(net117),
    .D(_0172_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfxtp_1 _6866_ (.CLK(net118),
    .D(_0173_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfxtp_1 _6867_ (.CLK(net119),
    .D(_0174_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfxtp_1 _6868_ (.CLK(net120),
    .D(_0175_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfxtp_1 _6869_ (.CLK(net121),
    .D(_0176_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_1 _6870_ (.CLK(net122),
    .D(_0177_),
    .Q(\egd_top.BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6871_ (.CLK(net123),
    .D(_0178_),
    .Q(\egd_top.BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6872_ (.CLK(net124),
    .D(_0179_),
    .Q(\egd_top.BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6873_ (.CLK(net125),
    .D(_0180_),
    .Q(\egd_top.BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6874_ (.CLK(net126),
    .D(_0181_),
    .Q(\egd_top.BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6875_ (.CLK(net127),
    .D(_0182_),
    .Q(\egd_top.BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6876_ (.CLK(net128),
    .D(_0183_),
    .Q(\egd_top.BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6877_ (.CLK(net129),
    .D(_0184_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfxtp_2 _6878_ (.CLK(net130),
    .D(_0185_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfxtp_2 _6879_ (.CLK(net131),
    .D(_0186_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfxtp_2 _6880_ (.CLK(net132),
    .D(_0187_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfxtp_1 _6881_ (.CLK(net133),
    .D(_0188_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfxtp_1 _6882_ (.CLK(net134),
    .D(_0189_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfxtp_1 _6883_ (.CLK(net135),
    .D(_0190_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfxtp_1 _6884_ (.CLK(net136),
    .D(_0191_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfxtp_1 _6885_ (.CLK(net137),
    .D(_0192_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfxtp_1 _6886_ (.CLK(net138),
    .D(_0193_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfxtp_1 _6887_ (.CLK(net139),
    .D(_0194_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfxtp_1 _6888_ (.CLK(net140),
    .D(_0195_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfxtp_1 _6889_ (.CLK(net141),
    .D(_0196_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfxtp_1 _6890_ (.CLK(net142),
    .D(_0197_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfxtp_1 _6891_ (.CLK(net143),
    .D(_0198_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfxtp_1 _6892_ (.CLK(net144),
    .D(_0199_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfxtp_1 _6893_ (.CLK(net145),
    .D(_0200_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfxtp_1 _6894_ (.CLK(net146),
    .D(_0201_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfxtp_1 _6895_ (.CLK(net147),
    .D(_0202_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfxtp_1 _6896_ (.CLK(net148),
    .D(_0203_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfxtp_1 _6897_ (.CLK(net149),
    .D(_0204_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfxtp_1 _6898_ (.CLK(net150),
    .D(_0205_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfxtp_1 _6899_ (.CLK(net151),
    .D(_0206_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _6900_ (.CLK(net152),
    .D(_0207_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _6901_ (.CLK(net153),
    .D(_0208_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(net154),
    .D(_0209_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _6903_ (.CLK(net155),
    .D(_0210_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _6904_ (.CLK(net156),
    .D(_0211_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _6905_ (.CLK(net157),
    .D(_0212_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(net158),
    .D(_0213_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(net159),
    .D(_0214_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(net160),
    .D(_0215_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _6909_ (.CLK(net161),
    .D(_0216_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _6910_ (.CLK(net162),
    .D(_0217_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _6911_ (.CLK(net163),
    .D(_0218_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _6912_ (.CLK(net164),
    .D(_0219_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _6913_ (.CLK(net165),
    .D(_0220_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _6914_ (.CLK(net166),
    .D(_0221_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _6915_ (.CLK(net167),
    .D(_0222_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _6916_ (.CLK(net168),
    .D(_0223_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _6917_ (.CLK(net169),
    .D(_0224_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _6918_ (.CLK(net170),
    .D(_0225_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _6919_ (.CLK(net171),
    .D(_0226_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _6920_ (.CLK(net172),
    .D(_0227_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _6921_ (.CLK(net173),
    .D(_0228_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _6922_ (.CLK(net174),
    .D(_0229_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _6923_ (.CLK(net175),
    .D(_0230_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _6924_ (.CLK(net176),
    .D(_0231_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _6925_ (.CLK(net177),
    .D(_0232_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _6926_ (.CLK(net178),
    .D(_0233_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _6927_ (.CLK(net179),
    .D(_0234_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _6928_ (.CLK(net180),
    .D(_0235_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _6929_ (.CLK(net181),
    .D(_0236_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _6930_ (.CLK(net182),
    .D(_0237_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _6931_ (.CLK(net183),
    .D(_0238_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _6932_ (.CLK(net184),
    .D(_0239_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _6933_ (.CLK(net185),
    .D(_0240_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _6934_ (.CLK(net186),
    .D(_0241_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _6935_ (.CLK(net187),
    .D(_0242_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _6936_ (.CLK(net188),
    .D(_0243_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _6937_ (.CLK(net189),
    .D(_0244_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _6938_ (.CLK(net190),
    .D(_0245_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _6939_ (.CLK(net191),
    .D(_0246_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _6940_ (.CLK(net192),
    .D(_0247_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6941_ (.CLK(net193),
    .D(_0248_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6942_ (.CLK(net194),
    .D(_0249_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6943_ (.CLK(net195),
    .D(_0250_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6944_ (.CLK(net36),
    .D(_0251_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6945_ (.CLK(net37),
    .D(_0252_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6946_ (.CLK(net38),
    .D(_0253_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6947_ (.CLK(net39),
    .D(_0254_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6948_ (.CLK(net40),
    .D(_0255_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6949_ (.CLK(net41),
    .D(_0256_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6950_ (.CLK(net42),
    .D(_0257_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6951_ (.CLK(net43),
    .D(_0258_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6952_ (.CLK(net44),
    .D(_0259_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6953_ (.CLK(net45),
    .D(_0260_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6954_ (.CLK(net46),
    .D(_0261_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6955_ (.CLK(net47),
    .D(_0262_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_2 _6956_ (.CLK(net48),
    .D(_0263_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _6957_ (.CLK(net49),
    .D(_0264_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_2 _6958_ (.CLK(net50),
    .D(_0265_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _6959_ (.CLK(net51),
    .D(_0266_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _6960_ (.CLK(net52),
    .D(_0267_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6961_ (.CLK(net53),
    .D(_0268_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _6962_ (.CLK(net54),
    .D(_0269_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6963_ (.CLK(net55),
    .D(_0270_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6964_ (.CLK(net56),
    .D(_0271_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _6965_ (.CLK(net57),
    .D(_0272_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6966_ (.CLK(net58),
    .D(_0273_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6967_ (.CLK(net59),
    .D(_0274_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6968_ (.CLK(net60),
    .D(_0275_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6969_ (.CLK(net61),
    .D(_0276_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6970_ (.CLK(net62),
    .D(_0277_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6971_ (.CLK(net63),
    .D(_0278_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6972_ (.CLK(net64),
    .D(_0279_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6973_ (.CLK(net65),
    .D(_0280_),
    .Q(\egd_top.BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6974_ (.CLK(net66),
    .D(_0281_),
    .Q(\egd_top.BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(net67),
    .D(_0282_),
    .Q(\egd_top.BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(net68),
    .D(_0283_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(net69),
    .D(_0284_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(net70),
    .D(_0285_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(net71),
    .D(_0286_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6980_ (.CLK(net72),
    .D(_0287_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(net73),
    .D(_0288_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6982_ (.CLK(net74),
    .D(_0289_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(net75),
    .D(_0290_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(net76),
    .D(_0291_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(net77),
    .D(_0292_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6986_ (.CLK(net78),
    .D(_0293_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(net79),
    .D(_0294_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6988_ (.CLK(net80),
    .D(_0295_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(net81),
    .D(_0296_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6990_ (.CLK(net82),
    .D(_0297_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6991_ (.CLK(net83),
    .D(_0298_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfxtp_1 _6992_ (.CLK(net84),
    .D(_0299_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfxtp_1 _6993_ (.CLK(net85),
    .D(_0300_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfxtp_1 _6994_ (.CLK(net86),
    .D(_0301_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfxtp_1 _6995_ (.CLK(net87),
    .D(_0302_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(net88),
    .D(_0303_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfxtp_1 _6997_ (.CLK(net89),
    .D(_0304_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfxtp_1 _6998_ (.CLK(net90),
    .D(_0305_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfxtp_1 _6999_ (.CLK(net91),
    .D(_0306_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfxtp_1 _7000_ (.CLK(net92),
    .D(_0307_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfxtp_1 _7001_ (.CLK(net93),
    .D(_0308_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfxtp_1 _7002_ (.CLK(net94),
    .D(_0309_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfxtp_1 _7003_ (.CLK(net95),
    .D(_0310_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfxtp_1 _7004_ (.CLK(net96),
    .D(_0311_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfxtp_1 _7005_ (.CLK(net97),
    .D(_0312_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfxtp_1 _7006_ (.CLK(net98),
    .D(_0313_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfxtp_1 _7007_ (.CLK(net99),
    .D(_0314_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfxtp_2 _7008_ (.CLK(net100),
    .D(_0315_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_2 _7009_ (.CLK(net101),
    .D(_0316_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _7010_ (.CLK(net102),
    .D(_0317_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _7011_ (.CLK(net103),
    .D(_0318_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_2 _7012_ (.CLK(net104),
    .D(_0319_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _7013_ (.CLK(net105),
    .D(_0320_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _7014_ (.CLK(net35),
    .D(_0321_),
    .Q(net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2958_ (.A(_2958_),
    .X(clknet_0__2958_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2959_ (.A(_2959_),
    .X(clknet_0__2959_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2960_ (.A(_2960_),
    .X(clknet_0__2960_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2961_ (.A(_2961_),
    .X(clknet_0__2961_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2962_ (.A(_2962_),
    .X(clknet_0__2962_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2963_ (.A(_2963_),
    .X(clknet_0__2963_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2964_ (.A(_2964_),
    .X(clknet_0__2964_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2965_ (.A(_2965_),
    .X(clknet_0__2965_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2966_ (.A(_2966_),
    .X(clknet_0__2966_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2967_ (.A(_2967_),
    .X(clknet_0__2967_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2968_ (.A(_2968_),
    .X(clknet_0__2968_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2969_ (.A(_2969_),
    .X(clknet_0__2969_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2970_ (.A(_2970_),
    .X(clknet_0__2970_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2971_ (.A(_2971_),
    .X(clknet_0__2971_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2972_ (.A(_2972_),
    .X(clknet_0__2972_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2973_ (.A(_2973_),
    .X(clknet_0__2973_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2974_ (.A(_2974_),
    .X(clknet_0__2974_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2975_ (.A(_2975_),
    .X(clknet_0__2975_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2958_ (.A(clknet_0__2958_),
    .X(clknet_1_0__leaf__2958_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2959_ (.A(clknet_0__2959_),
    .X(clknet_1_0__leaf__2959_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2960_ (.A(clknet_0__2960_),
    .X(clknet_1_0__leaf__2960_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2961_ (.A(clknet_0__2961_),
    .X(clknet_1_0__leaf__2961_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2962_ (.A(clknet_0__2962_),
    .X(clknet_1_0__leaf__2962_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2963_ (.A(clknet_0__2963_),
    .X(clknet_1_0__leaf__2963_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2964_ (.A(clknet_0__2964_),
    .X(clknet_1_0__leaf__2964_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2965_ (.A(clknet_0__2965_),
    .X(clknet_1_0__leaf__2965_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2966_ (.A(clknet_0__2966_),
    .X(clknet_1_0__leaf__2966_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2967_ (.A(clknet_0__2967_),
    .X(clknet_1_0__leaf__2967_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2968_ (.A(clknet_0__2968_),
    .X(clknet_1_0__leaf__2968_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2969_ (.A(clknet_0__2969_),
    .X(clknet_1_0__leaf__2969_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2970_ (.A(clknet_0__2970_),
    .X(clknet_1_0__leaf__2970_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2971_ (.A(clknet_0__2971_),
    .X(clknet_1_0__leaf__2971_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2972_ (.A(clknet_0__2972_),
    .X(clknet_1_0__leaf__2972_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2973_ (.A(clknet_0__2973_),
    .X(clknet_1_0__leaf__2973_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2974_ (.A(clknet_0__2974_),
    .X(clknet_1_0__leaf__2974_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2975_ (.A(clknet_0__2975_),
    .X(clknet_1_0__leaf__2975_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2958_ (.A(clknet_0__2958_),
    .X(clknet_1_1__leaf__2958_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2959_ (.A(clknet_0__2959_),
    .X(clknet_1_1__leaf__2959_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2960_ (.A(clknet_0__2960_),
    .X(clknet_1_1__leaf__2960_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2961_ (.A(clknet_0__2961_),
    .X(clknet_1_1__leaf__2961_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2962_ (.A(clknet_0__2962_),
    .X(clknet_1_1__leaf__2962_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2963_ (.A(clknet_0__2963_),
    .X(clknet_1_1__leaf__2963_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2964_ (.A(clknet_0__2964_),
    .X(clknet_1_1__leaf__2964_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2965_ (.A(clknet_0__2965_),
    .X(clknet_1_1__leaf__2965_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2966_ (.A(clknet_0__2966_),
    .X(clknet_1_1__leaf__2966_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2967_ (.A(clknet_0__2967_),
    .X(clknet_1_1__leaf__2967_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2968_ (.A(clknet_0__2968_),
    .X(clknet_1_1__leaf__2968_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2969_ (.A(clknet_0__2969_),
    .X(clknet_1_1__leaf__2969_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2970_ (.A(clknet_0__2970_),
    .X(clknet_1_1__leaf__2970_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2971_ (.A(clknet_0__2971_),
    .X(clknet_1_1__leaf__2971_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2972_ (.A(clknet_0__2972_),
    .X(clknet_1_1__leaf__2972_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2973_ (.A(clknet_0__2973_),
    .X(clknet_1_1__leaf__2973_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2974_ (.A(clknet_0__2974_),
    .X(clknet_1_1__leaf__2974_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2975_ (.A(clknet_0__2975_),
    .X(clknet_1_1__leaf__2975_));
 sky130_fd_sc_hd__buf_1 hold1 (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_3019_),
    .X(net197));
 sky130_fd_sc_hd__buf_1 hold3 (.A(\egd_top.BitStream_buffer.buffer_index[5] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_2450_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net29),
    .X(net202));
 sky130_fd_sc_hd__buf_4 input1 (.A(la_data_in_47_32[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(la_data_in_47_32[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(la_data_in_47_32[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(la_data_in_47_32[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(la_data_in_47_32[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(la_data_in_47_32[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(la_data_in_47_32[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(la_data_in_47_32[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(la_data_in_49_48[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(la_data_in_49_48[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(la_data_in_65),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(la_data_in_47_32[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(la_data_in_47_32[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(la_data_in_47_32[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(la_data_in_47_32[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(la_data_in_47_32[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(la_data_in_47_32[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(la_data_in_47_32[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(la_data_in_47_32[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(la_data_out_15_8[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(la_data_out_15_8[1]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(la_data_out_15_8[2]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(la_data_out_15_8[3]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(la_data_out_15_8[4]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(la_data_out_15_8[5]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(la_data_out_15_8[6]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_data_out_15_8[7]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(la_data_out_18_16[0]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(la_data_out_18_16[1]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(la_data_out_18_16[2]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(la_data_out_22_19[0]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(la_data_out_22_19[1]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(la_data_out_22_19[2]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(la_data_out_22_19[3]));
endmodule

