magic
tech sky130A
magscale 1 2
timestamp 1695970226
<< obsli1 >>
rect 1104 2159 49956 50609
<< obsm1 >>
rect 1104 1572 49956 50640
<< metal2 >>
rect 1214 0 1270 800
rect 2686 0 2742 800
rect 4158 0 4214 800
rect 5630 0 5686 800
rect 7102 0 7158 800
rect 8574 0 8630 800
rect 10046 0 10102 800
rect 11518 0 11574 800
rect 12990 0 13046 800
rect 14462 0 14518 800
rect 15934 0 15990 800
rect 17406 0 17462 800
rect 18878 0 18934 800
rect 20350 0 20406 800
rect 21822 0 21878 800
rect 23294 0 23350 800
rect 24766 0 24822 800
rect 26238 0 26294 800
rect 27710 0 27766 800
rect 29182 0 29238 800
rect 30654 0 30710 800
rect 32126 0 32182 800
rect 33598 0 33654 800
rect 35070 0 35126 800
rect 36542 0 36598 800
rect 38014 0 38070 800
rect 39486 0 39542 800
rect 40958 0 41014 800
rect 42430 0 42486 800
rect 43902 0 43958 800
rect 45374 0 45430 800
rect 46846 0 46902 800
rect 48318 0 48374 800
rect 49790 0 49846 800
<< obsm2 >>
rect 1216 856 49844 50629
rect 1326 734 2630 856
rect 2798 734 4102 856
rect 4270 734 5574 856
rect 5742 734 7046 856
rect 7214 734 8518 856
rect 8686 734 9990 856
rect 10158 734 11462 856
rect 11630 734 12934 856
rect 13102 734 14406 856
rect 14574 734 15878 856
rect 16046 734 17350 856
rect 17518 734 18822 856
rect 18990 734 20294 856
rect 20462 734 21766 856
rect 21934 734 23238 856
rect 23406 734 24710 856
rect 24878 734 26182 856
rect 26350 734 27654 856
rect 27822 734 29126 856
rect 29294 734 30598 856
rect 30766 734 32070 856
rect 32238 734 33542 856
rect 33710 734 35014 856
rect 35182 734 36486 856
rect 36654 734 37958 856
rect 38126 734 39430 856
rect 39598 734 40902 856
rect 41070 734 42374 856
rect 42542 734 43846 856
rect 44014 734 45318 856
rect 45486 734 46790 856
rect 46958 734 48262 856
rect 48430 734 49734 856
<< metal3 >>
rect 0 26392 800 26512
<< obsm3 >>
rect 800 26592 48379 50625
rect 880 26312 48379 26592
rect 800 1803 48379 26312
<< metal4 >>
rect 4208 2128 4528 50640
rect 19568 2128 19888 50640
rect 34928 2128 35248 50640
<< obsm4 >>
rect 12571 2048 19488 42533
rect 19968 2048 34848 42533
rect 35328 2048 46861 42533
rect 12571 1803 46861 2048
<< labels >>
rlabel metal2 s 23294 0 23350 800 6 la_data_in_47_32[0]
port 1 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in_47_32[10]
port 2 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in_47_32[11]
port 3 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in_47_32[12]
port 4 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 la_data_in_47_32[13]
port 5 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in_47_32[14]
port 6 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in_47_32[15]
port 7 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in_47_32[1]
port 8 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in_47_32[2]
port 9 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in_47_32[3]
port 10 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_data_in_47_32[4]
port 11 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in_47_32[5]
port 12 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_data_in_47_32[6]
port 13 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in_47_32[7]
port 14 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in_47_32[8]
port 15 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_data_in_47_32[9]
port 16 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in_49_48[0]
port 17 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in_49_48[1]
port 18 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in_65
port 19 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 la_data_out_15_8[0]
port 20 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 la_data_out_15_8[1]
port 21 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 la_data_out_15_8[2]
port 22 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 la_data_out_15_8[3]
port 23 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 la_data_out_15_8[4]
port 24 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 la_data_out_15_8[5]
port 25 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 la_data_out_15_8[6]
port 26 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 la_data_out_15_8[7]
port 27 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 la_data_out_18_16[0]
port 28 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 la_data_out_18_16[1]
port 29 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 la_data_out_18_16[2]
port 30 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out_22_19[0]
port 31 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 la_data_out_22_19[1]
port 32 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 la_data_out_22_19[2]
port 33 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 la_data_out_22_19[3]
port 34 nsew signal output
rlabel metal4 s 4208 2128 4528 50640 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 50640 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 50640 6 vssd1
port 36 nsew ground bidirectional
rlabel metal3 s 0 26392 800 26512 6 wb_clk_i
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 51094 53238
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9417636
string GDS_FILE /home/uniccass/H.264_Decoder/openlane/egd_top_wrapper/runs/23_09_28_23_25/results/signoff/egd_top_wrapper.magic.gds
string GDS_START 510854
<< end >>

