VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO egd_top_wrapper
  CLASS BLOCK ;
  FOREIGN egd_top_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 266.840 BY 277.560 ;
  PIN la_data_in_47_32[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END la_data_in_47_32[0]
  PIN la_data_in_47_32[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END la_data_in_47_32[10]
  PIN la_data_in_47_32[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END la_data_in_47_32[11]
  PIN la_data_in_47_32[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END la_data_in_47_32[12]
  PIN la_data_in_47_32[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END la_data_in_47_32[13]
  PIN la_data_in_47_32[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END la_data_in_47_32[14]
  PIN la_data_in_47_32[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END la_data_in_47_32[15]
  PIN la_data_in_47_32[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END la_data_in_47_32[1]
  PIN la_data_in_47_32[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END la_data_in_47_32[2]
  PIN la_data_in_47_32[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END la_data_in_47_32[3]
  PIN la_data_in_47_32[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END la_data_in_47_32[4]
  PIN la_data_in_47_32[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END la_data_in_47_32[5]
  PIN la_data_in_47_32[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END la_data_in_47_32[6]
  PIN la_data_in_47_32[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END la_data_in_47_32[7]
  PIN la_data_in_47_32[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END la_data_in_47_32[8]
  PIN la_data_in_47_32[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END la_data_in_47_32[9]
  PIN la_data_in_49_48[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END la_data_in_49_48[0]
  PIN la_data_in_49_48[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_data_in_49_48[1]
  PIN la_data_in_65
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_data_in_65
  PIN la_data_out_15_8[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END la_data_out_15_8[0]
  PIN la_data_out_15_8[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END la_data_out_15_8[1]
  PIN la_data_out_15_8[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END la_data_out_15_8[2]
  PIN la_data_out_15_8[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END la_data_out_15_8[3]
  PIN la_data_out_15_8[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END la_data_out_15_8[4]
  PIN la_data_out_15_8[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END la_data_out_15_8[5]
  PIN la_data_out_15_8[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END la_data_out_15_8[6]
  PIN la_data_out_15_8[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END la_data_out_15_8[7]
  PIN la_data_out_18_16[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END la_data_out_18_16[0]
  PIN la_data_out_18_16[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END la_data_out_18_16[1]
  PIN la_data_out_18_16[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END la_data_out_18_16[2]
  PIN la_data_out_22_19[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END la_data_out_22_19[0]
  PIN la_data_out_22_19[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END la_data_out_22_19[1]
  PIN la_data_out_22_19[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END la_data_out_22_19[2]
  PIN la_data_out_22_19[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END la_data_out_22_19[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 266.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 266.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 266.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 261.280 266.645 ;
      LAYER met1 ;
        RECT 4.210 9.220 266.730 266.800 ;
      LAYER met2 ;
        RECT 4.240 4.280 266.710 266.745 ;
        RECT 4.790 3.670 11.770 4.280 ;
        RECT 12.610 3.670 19.590 4.280 ;
        RECT 20.430 3.670 27.410 4.280 ;
        RECT 28.250 3.670 35.230 4.280 ;
        RECT 36.070 3.670 43.050 4.280 ;
        RECT 43.890 3.670 50.870 4.280 ;
        RECT 51.710 3.670 58.690 4.280 ;
        RECT 59.530 3.670 66.510 4.280 ;
        RECT 67.350 3.670 74.330 4.280 ;
        RECT 75.170 3.670 82.150 4.280 ;
        RECT 82.990 3.670 89.970 4.280 ;
        RECT 90.810 3.670 97.790 4.280 ;
        RECT 98.630 3.670 105.610 4.280 ;
        RECT 106.450 3.670 113.430 4.280 ;
        RECT 114.270 3.670 121.250 4.280 ;
        RECT 122.090 3.670 129.070 4.280 ;
        RECT 129.910 3.670 136.890 4.280 ;
        RECT 137.730 3.670 144.710 4.280 ;
        RECT 145.550 3.670 152.530 4.280 ;
        RECT 153.370 3.670 160.350 4.280 ;
        RECT 161.190 3.670 168.170 4.280 ;
        RECT 169.010 3.670 175.990 4.280 ;
        RECT 176.830 3.670 183.810 4.280 ;
        RECT 184.650 3.670 191.630 4.280 ;
        RECT 192.470 3.670 199.450 4.280 ;
        RECT 200.290 3.670 207.270 4.280 ;
        RECT 208.110 3.670 215.090 4.280 ;
        RECT 215.930 3.670 222.910 4.280 ;
        RECT 223.750 3.670 230.730 4.280 ;
        RECT 231.570 3.670 238.550 4.280 ;
        RECT 239.390 3.670 246.370 4.280 ;
        RECT 247.210 3.670 254.190 4.280 ;
        RECT 255.030 3.670 262.010 4.280 ;
        RECT 262.850 3.670 266.710 4.280 ;
      LAYER met3 ;
        RECT 4.000 138.400 266.735 266.725 ;
        RECT 4.400 137.000 266.735 138.400 ;
        RECT 4.000 10.715 266.735 137.000 ;
      LAYER met4 ;
        RECT 33.415 11.735 97.440 224.905 ;
        RECT 99.840 11.735 174.240 224.905 ;
        RECT 176.640 11.735 251.040 224.905 ;
        RECT 253.440 11.735 266.505 224.905 ;
  END
END egd_top_wrapper
END LIBRARY

