// This is the unpowered netlist.
module egd_top (clk,
    reset_n,
    BitStream_buffer_input,
    exp_golomb_decoding_output,
    exp_golomb_sel,
    half_fill_counter,
    reset_counter);
 input clk;
 input reset_n;
 input [15:0] BitStream_buffer_input;
 output [7:0] exp_golomb_decoding_output;
 input [1:0] exp_golomb_sel;
 output [2:0] half_fill_counter;
 output [3:0] reset_counter;

 wire \BitStream_buffer.BS_buffer[0] ;
 wire \BitStream_buffer.BS_buffer[100] ;
 wire \BitStream_buffer.BS_buffer[101] ;
 wire \BitStream_buffer.BS_buffer[102] ;
 wire \BitStream_buffer.BS_buffer[103] ;
 wire \BitStream_buffer.BS_buffer[104] ;
 wire \BitStream_buffer.BS_buffer[105] ;
 wire \BitStream_buffer.BS_buffer[106] ;
 wire \BitStream_buffer.BS_buffer[107] ;
 wire \BitStream_buffer.BS_buffer[108] ;
 wire \BitStream_buffer.BS_buffer[109] ;
 wire \BitStream_buffer.BS_buffer[10] ;
 wire \BitStream_buffer.BS_buffer[110] ;
 wire \BitStream_buffer.BS_buffer[111] ;
 wire \BitStream_buffer.BS_buffer[112] ;
 wire \BitStream_buffer.BS_buffer[113] ;
 wire \BitStream_buffer.BS_buffer[114] ;
 wire \BitStream_buffer.BS_buffer[115] ;
 wire \BitStream_buffer.BS_buffer[116] ;
 wire \BitStream_buffer.BS_buffer[117] ;
 wire \BitStream_buffer.BS_buffer[118] ;
 wire \BitStream_buffer.BS_buffer[119] ;
 wire \BitStream_buffer.BS_buffer[11] ;
 wire \BitStream_buffer.BS_buffer[120] ;
 wire \BitStream_buffer.BS_buffer[121] ;
 wire \BitStream_buffer.BS_buffer[122] ;
 wire \BitStream_buffer.BS_buffer[123] ;
 wire \BitStream_buffer.BS_buffer[124] ;
 wire \BitStream_buffer.BS_buffer[125] ;
 wire \BitStream_buffer.BS_buffer[126] ;
 wire \BitStream_buffer.BS_buffer[127] ;
 wire \BitStream_buffer.BS_buffer[12] ;
 wire \BitStream_buffer.BS_buffer[13] ;
 wire \BitStream_buffer.BS_buffer[14] ;
 wire \BitStream_buffer.BS_buffer[15] ;
 wire \BitStream_buffer.BS_buffer[16] ;
 wire \BitStream_buffer.BS_buffer[17] ;
 wire \BitStream_buffer.BS_buffer[18] ;
 wire \BitStream_buffer.BS_buffer[19] ;
 wire \BitStream_buffer.BS_buffer[1] ;
 wire \BitStream_buffer.BS_buffer[20] ;
 wire \BitStream_buffer.BS_buffer[21] ;
 wire \BitStream_buffer.BS_buffer[22] ;
 wire \BitStream_buffer.BS_buffer[23] ;
 wire \BitStream_buffer.BS_buffer[24] ;
 wire \BitStream_buffer.BS_buffer[25] ;
 wire \BitStream_buffer.BS_buffer[26] ;
 wire \BitStream_buffer.BS_buffer[27] ;
 wire \BitStream_buffer.BS_buffer[28] ;
 wire \BitStream_buffer.BS_buffer[29] ;
 wire \BitStream_buffer.BS_buffer[2] ;
 wire \BitStream_buffer.BS_buffer[30] ;
 wire \BitStream_buffer.BS_buffer[31] ;
 wire \BitStream_buffer.BS_buffer[32] ;
 wire \BitStream_buffer.BS_buffer[33] ;
 wire \BitStream_buffer.BS_buffer[34] ;
 wire \BitStream_buffer.BS_buffer[35] ;
 wire \BitStream_buffer.BS_buffer[36] ;
 wire \BitStream_buffer.BS_buffer[37] ;
 wire \BitStream_buffer.BS_buffer[38] ;
 wire \BitStream_buffer.BS_buffer[39] ;
 wire \BitStream_buffer.BS_buffer[3] ;
 wire \BitStream_buffer.BS_buffer[40] ;
 wire \BitStream_buffer.BS_buffer[41] ;
 wire \BitStream_buffer.BS_buffer[42] ;
 wire \BitStream_buffer.BS_buffer[43] ;
 wire \BitStream_buffer.BS_buffer[44] ;
 wire \BitStream_buffer.BS_buffer[45] ;
 wire \BitStream_buffer.BS_buffer[46] ;
 wire \BitStream_buffer.BS_buffer[47] ;
 wire \BitStream_buffer.BS_buffer[48] ;
 wire \BitStream_buffer.BS_buffer[49] ;
 wire \BitStream_buffer.BS_buffer[4] ;
 wire \BitStream_buffer.BS_buffer[50] ;
 wire \BitStream_buffer.BS_buffer[51] ;
 wire \BitStream_buffer.BS_buffer[52] ;
 wire \BitStream_buffer.BS_buffer[53] ;
 wire \BitStream_buffer.BS_buffer[54] ;
 wire \BitStream_buffer.BS_buffer[55] ;
 wire \BitStream_buffer.BS_buffer[56] ;
 wire \BitStream_buffer.BS_buffer[57] ;
 wire \BitStream_buffer.BS_buffer[58] ;
 wire \BitStream_buffer.BS_buffer[59] ;
 wire \BitStream_buffer.BS_buffer[5] ;
 wire \BitStream_buffer.BS_buffer[60] ;
 wire \BitStream_buffer.BS_buffer[61] ;
 wire \BitStream_buffer.BS_buffer[62] ;
 wire \BitStream_buffer.BS_buffer[63] ;
 wire \BitStream_buffer.BS_buffer[64] ;
 wire \BitStream_buffer.BS_buffer[65] ;
 wire \BitStream_buffer.BS_buffer[66] ;
 wire \BitStream_buffer.BS_buffer[67] ;
 wire \BitStream_buffer.BS_buffer[68] ;
 wire \BitStream_buffer.BS_buffer[69] ;
 wire \BitStream_buffer.BS_buffer[6] ;
 wire \BitStream_buffer.BS_buffer[70] ;
 wire \BitStream_buffer.BS_buffer[71] ;
 wire \BitStream_buffer.BS_buffer[72] ;
 wire \BitStream_buffer.BS_buffer[73] ;
 wire \BitStream_buffer.BS_buffer[74] ;
 wire \BitStream_buffer.BS_buffer[75] ;
 wire \BitStream_buffer.BS_buffer[76] ;
 wire \BitStream_buffer.BS_buffer[77] ;
 wire \BitStream_buffer.BS_buffer[78] ;
 wire \BitStream_buffer.BS_buffer[79] ;
 wire \BitStream_buffer.BS_buffer[7] ;
 wire \BitStream_buffer.BS_buffer[80] ;
 wire \BitStream_buffer.BS_buffer[81] ;
 wire \BitStream_buffer.BS_buffer[82] ;
 wire \BitStream_buffer.BS_buffer[83] ;
 wire \BitStream_buffer.BS_buffer[84] ;
 wire \BitStream_buffer.BS_buffer[85] ;
 wire \BitStream_buffer.BS_buffer[86] ;
 wire \BitStream_buffer.BS_buffer[87] ;
 wire \BitStream_buffer.BS_buffer[88] ;
 wire \BitStream_buffer.BS_buffer[89] ;
 wire \BitStream_buffer.BS_buffer[8] ;
 wire \BitStream_buffer.BS_buffer[90] ;
 wire \BitStream_buffer.BS_buffer[91] ;
 wire \BitStream_buffer.BS_buffer[92] ;
 wire \BitStream_buffer.BS_buffer[93] ;
 wire \BitStream_buffer.BS_buffer[94] ;
 wire \BitStream_buffer.BS_buffer[95] ;
 wire \BitStream_buffer.BS_buffer[96] ;
 wire \BitStream_buffer.BS_buffer[97] ;
 wire \BitStream_buffer.BS_buffer[98] ;
 wire \BitStream_buffer.BS_buffer[99] ;
 wire \BitStream_buffer.BS_buffer[9] ;
 wire \BitStream_buffer.BitStream_buffer_output[10] ;
 wire \BitStream_buffer.BitStream_buffer_output[11] ;
 wire \BitStream_buffer.BitStream_buffer_output[12] ;
 wire \BitStream_buffer.BitStream_buffer_output[13] ;
 wire \BitStream_buffer.BitStream_buffer_output[14] ;
 wire \BitStream_buffer.BitStream_buffer_output[15] ;
 wire \BitStream_buffer.BitStream_buffer_output[1] ;
 wire \BitStream_buffer.BitStream_buffer_output[2] ;
 wire \BitStream_buffer.BitStream_buffer_output[3] ;
 wire \BitStream_buffer.BitStream_buffer_output[4] ;
 wire \BitStream_buffer.BitStream_buffer_output[5] ;
 wire \BitStream_buffer.BitStream_buffer_output[6] ;
 wire \BitStream_buffer.BitStream_buffer_output[7] ;
 wire \BitStream_buffer.BitStream_buffer_output[8] ;
 wire \BitStream_buffer.BitStream_buffer_output[9] ;
 wire \BitStream_buffer.BitStream_buffer_valid_n ;
 wire \BitStream_buffer.buffer_index[4] ;
 wire \BitStream_buffer.buffer_index[5] ;
 wire \BitStream_buffer.buffer_index[6] ;
 wire \BitStream_buffer.exp_golomb_len[1] ;
 wire \BitStream_buffer.exp_golomb_len[2] ;
 wire \BitStream_buffer.exp_golomb_len[3] ;
 wire \BitStream_buffer.pc[1] ;
 wire \BitStream_buffer.pc[2] ;
 wire \BitStream_buffer.pc[3] ;
 wire \BitStream_buffer.pc[4] ;
 wire \BitStream_buffer.pc[5] ;
 wire \BitStream_buffer.pc[6] ;
 wire \BitStream_buffer.pc_previous[0] ;
 wire \BitStream_buffer.pc_previous[1] ;
 wire \BitStream_buffer.pc_previous[2] ;
 wire \BitStream_buffer.pc_previous[3] ;
 wire \BitStream_buffer.pc_previous[4] ;
 wire \BitStream_buffer.pc_previous[5] ;
 wire \BitStream_buffer.pc_previous[6] ;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire clknet_0__2580_;
 wire clknet_0__2581_;
 wire clknet_0__2582_;
 wire clknet_0__2583_;
 wire clknet_0__2584_;
 wire clknet_0__2585_;
 wire clknet_0__2586_;
 wire clknet_0__2587_;
 wire clknet_0__2588_;
 wire clknet_0__2589_;
 wire clknet_0__2590_;
 wire clknet_0__2591_;
 wire clknet_0__2592_;
 wire clknet_0__2593_;
 wire clknet_0__2594_;
 wire clknet_0__2595_;
 wire clknet_0__2596_;
 wire clknet_0__2597_;
 wire clknet_1_0__leaf__2580_;
 wire clknet_1_0__leaf__2581_;
 wire clknet_1_0__leaf__2582_;
 wire clknet_1_0__leaf__2583_;
 wire clknet_1_0__leaf__2584_;
 wire clknet_1_0__leaf__2585_;
 wire clknet_1_0__leaf__2586_;
 wire clknet_1_0__leaf__2587_;
 wire clknet_1_0__leaf__2588_;
 wire clknet_1_0__leaf__2589_;
 wire clknet_1_0__leaf__2590_;
 wire clknet_1_0__leaf__2591_;
 wire clknet_1_0__leaf__2592_;
 wire clknet_1_0__leaf__2593_;
 wire clknet_1_0__leaf__2594_;
 wire clknet_1_0__leaf__2595_;
 wire clknet_1_0__leaf__2596_;
 wire clknet_1_0__leaf__2597_;
 wire clknet_1_1__leaf__2580_;
 wire clknet_1_1__leaf__2581_;
 wire clknet_1_1__leaf__2582_;
 wire clknet_1_1__leaf__2583_;
 wire clknet_1_1__leaf__2584_;
 wire clknet_1_1__leaf__2585_;
 wire clknet_1_1__leaf__2586_;
 wire clknet_1_1__leaf__2587_;
 wire clknet_1_1__leaf__2588_;
 wire clknet_1_1__leaf__2589_;
 wire clknet_1_1__leaf__2590_;
 wire clknet_1_1__leaf__2591_;
 wire clknet_1_1__leaf__2592_;
 wire clknet_1_1__leaf__2593_;
 wire clknet_1_1__leaf__2594_;
 wire clknet_1_1__leaf__2595_;
 wire clknet_1_1__leaf__2596_;
 wire clknet_1_1__leaf__2597_;
 wire \exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net13));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__buf_2 _3064_ (.A(\BitStream_buffer.BitStream_buffer_valid_n ),
    .X(_2598_));
 sky130_fd_sc_hd__buf_2 _3065_ (.A(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__inv_2 _3066_ (.A(\BitStream_buffer.pc[4] ),
    .Y(_2600_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(\BitStream_buffer.pc[5] ),
    .Y(_2601_));
 sky130_fd_sc_hd__and3_1 _3068_ (.A(_2600_),
    .B(_2601_),
    .C(\BitStream_buffer.pc[6] ),
    .X(_2602_));
 sky130_fd_sc_hd__inv_2 _3069_ (.A(_2602_),
    .Y(_2603_));
 sky130_fd_sc_hd__inv_2 _3070_ (.A(\BitStream_buffer.pc[3] ),
    .Y(_2604_));
 sky130_fd_sc_hd__inv_2 _3071_ (.A(net18),
    .Y(_2605_));
 sky130_fd_sc_hd__inv_2 _3072_ (.A(net17),
    .Y(_2606_));
 sky130_fd_sc_hd__nand2_4 _3073_ (.A(_2605_),
    .B(_2606_),
    .Y(_2607_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(_2607_),
    .Y(_2608_));
 sky130_fd_sc_hd__inv_2 _3075_ (.A(\BitStream_buffer.pc_previous[0] ),
    .Y(_2609_));
 sky130_fd_sc_hd__nand2_1 _3076_ (.A(_2608_),
    .B(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__nand2_4 _3077_ (.A(_2607_),
    .B(\BitStream_buffer.pc_previous[0] ),
    .Y(_2611_));
 sky130_fd_sc_hd__nand2_2 _3078_ (.A(_2610_),
    .B(_2611_),
    .Y(_2612_));
 sky130_fd_sc_hd__nand2_1 _3079_ (.A(_2612_),
    .B(\BitStream_buffer.pc[1] ),
    .Y(_2613_));
 sky130_fd_sc_hd__or3_1 _3080_ (.A(\BitStream_buffer.pc[2] ),
    .B(_2604_),
    .C(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__clkbuf_4 _3081_ (.A(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__nor2_2 _3082_ (.A(_2603_),
    .B(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__clkbuf_4 _3083_ (.A(_2616_),
    .X(_2617_));
 sky130_fd_sc_hd__inv_2 _3084_ (.A(_2612_),
    .Y(_2618_));
 sky130_fd_sc_hd__nand2_4 _3085_ (.A(_2618_),
    .B(\BitStream_buffer.pc[1] ),
    .Y(_2619_));
 sky130_fd_sc_hd__nor3_4 _3086_ (.A(\BitStream_buffer.pc[2] ),
    .B(_2604_),
    .C(_2619_),
    .Y(_2620_));
 sky130_fd_sc_hd__clkbuf_4 _3087_ (.A(_2602_),
    .X(_2621_));
 sky130_fd_sc_hd__and2_1 _3088_ (.A(_2620_),
    .B(_2621_),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_2 _3089_ (.A(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__clkbuf_4 _3090_ (.A(_2623_),
    .X(_2624_));
 sky130_fd_sc_hd__inv_2 _3091_ (.A(\BitStream_buffer.BS_buffer[73] ),
    .Y(_2625_));
 sky130_fd_sc_hd__inv_2 _3092_ (.A(\BitStream_buffer.pc[1] ),
    .Y(_2626_));
 sky130_fd_sc_hd__nand2_4 _3093_ (.A(_2618_),
    .B(_2626_),
    .Y(_2627_));
 sky130_fd_sc_hd__nor3_2 _3094_ (.A(\BitStream_buffer.pc[2] ),
    .B(_2604_),
    .C(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__nand2_2 _3095_ (.A(net35),
    .B(_2621_),
    .Y(_2629_));
 sky130_fd_sc_hd__clkbuf_4 _3096_ (.A(_2629_),
    .X(_2630_));
 sky130_fd_sc_hd__inv_2 _3097_ (.A(\BitStream_buffer.BS_buffer[72] ),
    .Y(_2631_));
 sky130_fd_sc_hd__nand2_1 _3098_ (.A(_2612_),
    .B(_2626_),
    .Y(_2632_));
 sky130_fd_sc_hd__or3_1 _3099_ (.A(\BitStream_buffer.pc[2] ),
    .B(_2604_),
    .C(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__buf_4 _3100_ (.A(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__or2_1 _3101_ (.A(_2603_),
    .B(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__clkbuf_2 _3102_ (.A(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__buf_6 _3103_ (.A(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__o22ai_1 _3104_ (.A1(_2625_),
    .A2(_2630_),
    .B1(_2631_),
    .B2(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__a221oi_1 _3105_ (.A1(\BitStream_buffer.BS_buffer[74] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[75] ),
    .B2(_2624_),
    .C1(_2638_),
    .Y(_2639_));
 sky130_fd_sc_hd__inv_2 _3106_ (.A(\BitStream_buffer.BS_buffer[64] ),
    .Y(_2640_));
 sky130_fd_sc_hd__inv_2 _3107_ (.A(_2632_),
    .Y(_2641_));
 sky130_fd_sc_hd__nor2_2 _3108_ (.A(\BitStream_buffer.pc[2] ),
    .B(\BitStream_buffer.pc[3] ),
    .Y(_2642_));
 sky130_fd_sc_hd__nand2_4 _3109_ (.A(_2641_),
    .B(_2642_),
    .Y(_2643_));
 sky130_fd_sc_hd__inv_2 _3110_ (.A(_2643_),
    .Y(_2644_));
 sky130_fd_sc_hd__nand2_2 _3111_ (.A(_2644_),
    .B(_2621_),
    .Y(_2645_));
 sky130_fd_sc_hd__clkbuf_4 _3112_ (.A(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__inv_2 _3113_ (.A(_2613_),
    .Y(_2647_));
 sky130_fd_sc_hd__nand2_4 _3114_ (.A(_2647_),
    .B(_2642_),
    .Y(_2648_));
 sky130_fd_sc_hd__nor2_2 _3115_ (.A(_2603_),
    .B(_2648_),
    .Y(_2649_));
 sky130_fd_sc_hd__buf_2 _3116_ (.A(_2649_),
    .X(_2650_));
 sky130_fd_sc_hd__nand2_1 _3117_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[66] ),
    .Y(_2651_));
 sky130_fd_sc_hd__inv_2 _3118_ (.A(\BitStream_buffer.BS_buffer[65] ),
    .Y(_2652_));
 sky130_fd_sc_hd__inv_2 _3119_ (.A(_2642_),
    .Y(_2653_));
 sky130_fd_sc_hd__nor2_4 _3120_ (.A(_2653_),
    .B(_2627_),
    .Y(_2654_));
 sky130_fd_sc_hd__nand2_1 _3121_ (.A(_2654_),
    .B(_2621_),
    .Y(_2655_));
 sky130_fd_sc_hd__clkbuf_2 _3122_ (.A(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__or2_1 _3123_ (.A(_2652_),
    .B(_2656_),
    .X(_2657_));
 sky130_fd_sc_hd__inv_2 _3124_ (.A(\BitStream_buffer.BS_buffer[67] ),
    .Y(_2658_));
 sky130_fd_sc_hd__nor2_4 _3125_ (.A(_2653_),
    .B(_2619_),
    .Y(_2659_));
 sky130_fd_sc_hd__nand2_1 _3126_ (.A(_2659_),
    .B(_2621_),
    .Y(_2660_));
 sky130_fd_sc_hd__clkbuf_2 _3127_ (.A(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__or2_1 _3128_ (.A(_2658_),
    .B(_2661_),
    .X(_2662_));
 sky130_fd_sc_hd__o2111a_1 _3129_ (.A1(_2640_),
    .A2(_2646_),
    .B1(_2651_),
    .C1(_2657_),
    .D1(_2662_),
    .X(_2663_));
 sky130_fd_sc_hd__inv_2 _3130_ (.A(\BitStream_buffer.BS_buffer[69] ),
    .Y(_2664_));
 sky130_fd_sc_hd__inv_2 _3131_ (.A(\BitStream_buffer.pc[2] ),
    .Y(_2665_));
 sky130_fd_sc_hd__nor2_2 _3132_ (.A(\BitStream_buffer.pc[3] ),
    .B(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__inv_2 _3133_ (.A(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__nor2_4 _3134_ (.A(_2667_),
    .B(_2627_),
    .Y(_2668_));
 sky130_fd_sc_hd__nand2_2 _3135_ (.A(_2668_),
    .B(_2621_),
    .Y(_2669_));
 sky130_fd_sc_hd__clkbuf_4 _3136_ (.A(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__inv_2 _3137_ (.A(\BitStream_buffer.BS_buffer[68] ),
    .Y(_2671_));
 sky130_fd_sc_hd__nand2_4 _3138_ (.A(_2641_),
    .B(_2666_),
    .Y(_2672_));
 sky130_fd_sc_hd__inv_2 _3139_ (.A(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__nand2_2 _3140_ (.A(_2673_),
    .B(_2621_),
    .Y(_2674_));
 sky130_fd_sc_hd__clkbuf_4 _3141_ (.A(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__o22ai_1 _3142_ (.A1(_2664_),
    .A2(_2670_),
    .B1(_2671_),
    .B2(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__nand2_4 _3143_ (.A(_2647_),
    .B(_2666_),
    .Y(_2677_));
 sky130_fd_sc_hd__nor2_2 _3144_ (.A(_2603_),
    .B(_2677_),
    .Y(_2678_));
 sky130_fd_sc_hd__clkbuf_4 _3145_ (.A(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__nor2_4 _3146_ (.A(_2667_),
    .B(_2619_),
    .Y(_2680_));
 sky130_fd_sc_hd__and2_2 _3147_ (.A(_2680_),
    .B(_2621_),
    .X(_2681_));
 sky130_fd_sc_hd__clkbuf_4 _3148_ (.A(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__a22o_1 _3149_ (.A1(\BitStream_buffer.BS_buffer[70] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[71] ),
    .X(_2683_));
 sky130_fd_sc_hd__nor2_1 _3150_ (.A(_2676_),
    .B(_2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__nand2_2 _3151_ (.A(\BitStream_buffer.pc[2] ),
    .B(\BitStream_buffer.pc[3] ),
    .Y(_2685_));
 sky130_fd_sc_hd__inv_2 _3152_ (.A(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__nand2_4 _3153_ (.A(_2647_),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__nor2_2 _3154_ (.A(_2603_),
    .B(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__buf_2 _3155_ (.A(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__nor2_4 _3156_ (.A(_2685_),
    .B(_2619_),
    .Y(_2690_));
 sky130_fd_sc_hd__and2_1 _3157_ (.A(_2690_),
    .B(_2602_),
    .X(_2691_));
 sky130_fd_sc_hd__clkbuf_2 _3158_ (.A(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__buf_2 _3159_ (.A(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__inv_2 _3160_ (.A(\BitStream_buffer.BS_buffer[77] ),
    .Y(_2694_));
 sky130_fd_sc_hd__nor2_4 _3161_ (.A(_2685_),
    .B(_2627_),
    .Y(_2695_));
 sky130_fd_sc_hd__nand2_2 _3162_ (.A(_2695_),
    .B(_2621_),
    .Y(_2696_));
 sky130_fd_sc_hd__clkbuf_4 _3163_ (.A(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__inv_2 _3164_ (.A(\BitStream_buffer.BS_buffer[76] ),
    .Y(_2698_));
 sky130_fd_sc_hd__nand2_4 _3165_ (.A(_2641_),
    .B(_2686_),
    .Y(_2699_));
 sky130_fd_sc_hd__inv_2 _3166_ (.A(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__nand2_2 _3167_ (.A(_2700_),
    .B(_2621_),
    .Y(_2701_));
 sky130_fd_sc_hd__buf_2 _3168_ (.A(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__o22ai_1 _3169_ (.A1(_2694_),
    .A2(_2697_),
    .B1(_2698_),
    .B2(_2702_),
    .Y(_2703_));
 sky130_fd_sc_hd__a221oi_1 _3170_ (.A1(\BitStream_buffer.BS_buffer[78] ),
    .A2(_2689_),
    .B1(\BitStream_buffer.BS_buffer[79] ),
    .B2(_2693_),
    .C1(_2703_),
    .Y(_2704_));
 sky130_fd_sc_hd__and4_1 _3171_ (.A(_2639_),
    .B(_2663_),
    .C(_2684_),
    .D(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__clkbuf_4 _3172_ (.A(\BitStream_buffer.BS_buffer[89] ),
    .X(_2706_));
 sky130_fd_sc_hd__inv_2 _3173_ (.A(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__inv_2 _3174_ (.A(\BitStream_buffer.pc[6] ),
    .Y(_2708_));
 sky130_fd_sc_hd__or3_1 _3175_ (.A(\BitStream_buffer.pc[5] ),
    .B(_2708_),
    .C(_2600_),
    .X(_2709_));
 sky130_fd_sc_hd__clkbuf_4 _3176_ (.A(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__inv_2 _3177_ (.A(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand2_2 _3178_ (.A(net35),
    .B(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__buf_2 _3179_ (.A(_2712_),
    .X(_2713_));
 sky130_fd_sc_hd__clkbuf_4 _3180_ (.A(\BitStream_buffer.BS_buffer[91] ),
    .X(_2714_));
 sky130_fd_sc_hd__inv_2 _3181_ (.A(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__nand2_2 _3182_ (.A(_2620_),
    .B(_2711_),
    .Y(_2716_));
 sky130_fd_sc_hd__clkbuf_2 _3183_ (.A(_2716_),
    .X(_2717_));
 sky130_fd_sc_hd__or2_1 _3184_ (.A(_2715_),
    .B(_2717_),
    .X(_2718_));
 sky130_fd_sc_hd__nor2_2 _3185_ (.A(_2710_),
    .B(_2615_),
    .Y(_2719_));
 sky130_fd_sc_hd__buf_4 _3186_ (.A(_2719_),
    .X(_2720_));
 sky130_fd_sc_hd__clkbuf_4 _3187_ (.A(\BitStream_buffer.BS_buffer[90] ),
    .X(_2721_));
 sky130_fd_sc_hd__nand2_1 _3188_ (.A(_2720_),
    .B(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__nor2_2 _3189_ (.A(_2710_),
    .B(_2634_),
    .Y(_2723_));
 sky130_fd_sc_hd__buf_4 _3190_ (.A(_2723_),
    .X(_2724_));
 sky130_fd_sc_hd__buf_2 _3191_ (.A(\BitStream_buffer.BS_buffer[88] ),
    .X(_2725_));
 sky130_fd_sc_hd__nand2_1 _3192_ (.A(_2724_),
    .B(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__o2111a_1 _3193_ (.A1(_2707_),
    .A2(_2713_),
    .B1(_2718_),
    .C1(_2722_),
    .D1(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__nor2_2 _3194_ (.A(_2710_),
    .B(_2687_),
    .Y(_2728_));
 sky130_fd_sc_hd__buf_2 _3195_ (.A(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__and2_1 _3196_ (.A(_2690_),
    .B(_2711_),
    .X(_2730_));
 sky130_fd_sc_hd__clkbuf_2 _3197_ (.A(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__buf_2 _3198_ (.A(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__inv_2 _3199_ (.A(\BitStream_buffer.BS_buffer[93] ),
    .Y(_2733_));
 sky130_fd_sc_hd__nand2_2 _3200_ (.A(_2695_),
    .B(_2711_),
    .Y(_2734_));
 sky130_fd_sc_hd__buf_2 _3201_ (.A(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__clkbuf_4 _3202_ (.A(\BitStream_buffer.BS_buffer[92] ),
    .X(_2736_));
 sky130_fd_sc_hd__inv_2 _3203_ (.A(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand2_2 _3204_ (.A(_2700_),
    .B(_2711_),
    .Y(_2738_));
 sky130_fd_sc_hd__buf_2 _3205_ (.A(_2738_),
    .X(_2739_));
 sky130_fd_sc_hd__o22ai_1 _3206_ (.A1(_2733_),
    .A2(_2735_),
    .B1(_2737_),
    .B2(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__a221oi_1 _3207_ (.A1(\BitStream_buffer.BS_buffer[94] ),
    .A2(_2729_),
    .B1(\BitStream_buffer.BS_buffer[95] ),
    .B2(_2732_),
    .C1(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__inv_2 _3208_ (.A(\BitStream_buffer.BS_buffer[81] ),
    .Y(_2742_));
 sky130_fd_sc_hd__nand2_2 _3209_ (.A(_2654_),
    .B(_2711_),
    .Y(_2743_));
 sky130_fd_sc_hd__buf_2 _3210_ (.A(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__nor2_2 _3211_ (.A(_2710_),
    .B(_2648_),
    .Y(_2745_));
 sky130_fd_sc_hd__buf_2 _3212_ (.A(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__nand2_1 _3213_ (.A(_2746_),
    .B(\BitStream_buffer.BS_buffer[82] ),
    .Y(_2747_));
 sky130_fd_sc_hd__nor2_2 _3214_ (.A(_2710_),
    .B(_2643_),
    .Y(_2748_));
 sky130_fd_sc_hd__buf_2 _3215_ (.A(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__nand2_1 _3216_ (.A(_2749_),
    .B(\BitStream_buffer.BS_buffer[80] ),
    .Y(_2750_));
 sky130_fd_sc_hd__inv_2 _3217_ (.A(\BitStream_buffer.BS_buffer[83] ),
    .Y(_2751_));
 sky130_fd_sc_hd__nand2_1 _3218_ (.A(_2659_),
    .B(_2711_),
    .Y(_2752_));
 sky130_fd_sc_hd__clkbuf_2 _3219_ (.A(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__or2_1 _3220_ (.A(_2751_),
    .B(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__o2111a_1 _3221_ (.A1(_2742_),
    .A2(_2744_),
    .B1(_2747_),
    .C1(_2750_),
    .D1(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__clkbuf_4 _3222_ (.A(\BitStream_buffer.BS_buffer[87] ),
    .X(_2756_));
 sky130_fd_sc_hd__inv_2 _3223_ (.A(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__nand2_2 _3224_ (.A(_2680_),
    .B(_2711_),
    .Y(_2758_));
 sky130_fd_sc_hd__buf_2 _3225_ (.A(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__nor2_2 _3226_ (.A(_2710_),
    .B(_2677_),
    .Y(_2760_));
 sky130_fd_sc_hd__buf_2 _3227_ (.A(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__clkbuf_4 _3228_ (.A(\BitStream_buffer.BS_buffer[86] ),
    .X(_2762_));
 sky130_fd_sc_hd__nand2_1 _3229_ (.A(_2761_),
    .B(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__nor2_2 _3230_ (.A(_2710_),
    .B(_2672_),
    .Y(_2764_));
 sky130_fd_sc_hd__buf_2 _3231_ (.A(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__buf_2 _3232_ (.A(\BitStream_buffer.BS_buffer[84] ),
    .X(_2766_));
 sky130_fd_sc_hd__nand2_1 _3233_ (.A(_2765_),
    .B(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__clkbuf_4 _3234_ (.A(\BitStream_buffer.BS_buffer[85] ),
    .X(_2768_));
 sky130_fd_sc_hd__inv_2 _3235_ (.A(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__nand2_1 _3236_ (.A(_2668_),
    .B(_2711_),
    .Y(_2770_));
 sky130_fd_sc_hd__clkbuf_2 _3237_ (.A(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__or2_1 _3238_ (.A(_2769_),
    .B(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__o2111a_1 _3239_ (.A1(_2757_),
    .A2(_2759_),
    .B1(_2763_),
    .C1(_2767_),
    .D1(_2772_),
    .X(_2773_));
 sky130_fd_sc_hd__and4_1 _3240_ (.A(_2727_),
    .B(_2741_),
    .C(_2755_),
    .D(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__inv_2 _3241_ (.A(\BitStream_buffer.BS_buffer[105] ),
    .Y(_2775_));
 sky130_fd_sc_hd__or3_1 _3242_ (.A(\BitStream_buffer.pc[4] ),
    .B(_2708_),
    .C(_2601_),
    .X(_2776_));
 sky130_fd_sc_hd__clkbuf_4 _3243_ (.A(_2776_),
    .X(_2777_));
 sky130_fd_sc_hd__inv_2 _3244_ (.A(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__nand2_2 _3245_ (.A(net35),
    .B(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__clkbuf_4 _3246_ (.A(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__clkbuf_4 _3247_ (.A(\BitStream_buffer.BS_buffer[107] ),
    .X(_2781_));
 sky130_fd_sc_hd__inv_2 _3248_ (.A(_2781_),
    .Y(_2782_));
 sky130_fd_sc_hd__nand2_1 _3249_ (.A(_2620_),
    .B(_2778_),
    .Y(_2783_));
 sky130_fd_sc_hd__clkbuf_2 _3250_ (.A(_2783_),
    .X(_2784_));
 sky130_fd_sc_hd__or2_1 _3251_ (.A(_2782_),
    .B(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__nor2_2 _3252_ (.A(_2777_),
    .B(_2615_),
    .Y(_2786_));
 sky130_fd_sc_hd__buf_4 _3253_ (.A(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__clkbuf_4 _3254_ (.A(\BitStream_buffer.BS_buffer[106] ),
    .X(_2788_));
 sky130_fd_sc_hd__nand2_1 _3255_ (.A(_2787_),
    .B(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__nor2_2 _3256_ (.A(_2777_),
    .B(_2634_),
    .Y(_2790_));
 sky130_fd_sc_hd__buf_4 _3257_ (.A(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__clkbuf_4 _3258_ (.A(\BitStream_buffer.BS_buffer[104] ),
    .X(_2792_));
 sky130_fd_sc_hd__nand2_1 _3259_ (.A(_2791_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__o2111a_1 _3260_ (.A1(_2775_),
    .A2(_2780_),
    .B1(_2785_),
    .C1(_2789_),
    .D1(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__inv_2 _3261_ (.A(\BitStream_buffer.BS_buffer[99] ),
    .Y(_2795_));
 sky130_fd_sc_hd__nand2_2 _3262_ (.A(_2659_),
    .B(_2778_),
    .Y(_2796_));
 sky130_fd_sc_hd__buf_2 _3263_ (.A(_2796_),
    .X(_2797_));
 sky130_fd_sc_hd__nor2_2 _3264_ (.A(_2777_),
    .B(_2643_),
    .Y(_2798_));
 sky130_fd_sc_hd__buf_2 _3265_ (.A(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__clkbuf_4 _3266_ (.A(\BitStream_buffer.BS_buffer[96] ),
    .X(_2800_));
 sky130_fd_sc_hd__nand2_1 _3267_ (.A(_2799_),
    .B(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__nor2_2 _3268_ (.A(_2777_),
    .B(_2648_),
    .Y(_2802_));
 sky130_fd_sc_hd__clkbuf_4 _3269_ (.A(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__clkbuf_4 _3270_ (.A(\BitStream_buffer.BS_buffer[98] ),
    .X(_2804_));
 sky130_fd_sc_hd__nand2_1 _3271_ (.A(_2803_),
    .B(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__inv_2 _3272_ (.A(\BitStream_buffer.BS_buffer[97] ),
    .Y(_2806_));
 sky130_fd_sc_hd__nand2_2 _3273_ (.A(_2654_),
    .B(_2778_),
    .Y(_2807_));
 sky130_fd_sc_hd__clkbuf_2 _3274_ (.A(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__or2_1 _3275_ (.A(_2806_),
    .B(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__o2111a_1 _3276_ (.A1(_2795_),
    .A2(_2797_),
    .B1(_2801_),
    .C1(_2805_),
    .D1(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__inv_2 _3277_ (.A(\BitStream_buffer.BS_buffer[103] ),
    .Y(_2811_));
 sky130_fd_sc_hd__nand2_2 _3278_ (.A(_2680_),
    .B(_2778_),
    .Y(_2812_));
 sky130_fd_sc_hd__buf_2 _3279_ (.A(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__nor2_2 _3280_ (.A(_2777_),
    .B(_2677_),
    .Y(_2814_));
 sky130_fd_sc_hd__buf_2 _3281_ (.A(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__clkbuf_4 _3282_ (.A(\BitStream_buffer.BS_buffer[102] ),
    .X(_2816_));
 sky130_fd_sc_hd__nand2_1 _3283_ (.A(_2815_),
    .B(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__nor2_2 _3284_ (.A(_2777_),
    .B(_2672_),
    .Y(_2818_));
 sky130_fd_sc_hd__clkbuf_4 _3285_ (.A(_2818_),
    .X(_2819_));
 sky130_fd_sc_hd__clkbuf_4 _3286_ (.A(\BitStream_buffer.BS_buffer[100] ),
    .X(_2820_));
 sky130_fd_sc_hd__nand2_1 _3287_ (.A(_2819_),
    .B(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__inv_2 _3288_ (.A(\BitStream_buffer.BS_buffer[101] ),
    .Y(_2822_));
 sky130_fd_sc_hd__nand2_1 _3289_ (.A(_2668_),
    .B(_2778_),
    .Y(_2823_));
 sky130_fd_sc_hd__clkbuf_2 _3290_ (.A(_2823_),
    .X(_2824_));
 sky130_fd_sc_hd__or2_1 _3291_ (.A(_2822_),
    .B(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__o2111a_1 _3292_ (.A1(_2811_),
    .A2(_2813_),
    .B1(_2817_),
    .C1(_2821_),
    .D1(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__inv_2 _3293_ (.A(\BitStream_buffer.BS_buffer[111] ),
    .Y(_2827_));
 sky130_fd_sc_hd__nand2_2 _3294_ (.A(_2690_),
    .B(_2778_),
    .Y(_2828_));
 sky130_fd_sc_hd__buf_2 _3295_ (.A(_2828_),
    .X(_2829_));
 sky130_fd_sc_hd__nor2_2 _3296_ (.A(_2777_),
    .B(_2699_),
    .Y(_2830_));
 sky130_fd_sc_hd__buf_2 _3297_ (.A(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__clkbuf_4 _3298_ (.A(\BitStream_buffer.BS_buffer[108] ),
    .X(_2832_));
 sky130_fd_sc_hd__nand2_1 _3299_ (.A(_2831_),
    .B(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__nor2_2 _3300_ (.A(_2777_),
    .B(_2687_),
    .Y(_2834_));
 sky130_fd_sc_hd__buf_2 _3301_ (.A(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__clkbuf_4 _3302_ (.A(\BitStream_buffer.BS_buffer[110] ),
    .X(_2836_));
 sky130_fd_sc_hd__nand2_1 _3303_ (.A(_2835_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__clkbuf_4 _3304_ (.A(\BitStream_buffer.BS_buffer[109] ),
    .X(_2838_));
 sky130_fd_sc_hd__inv_2 _3305_ (.A(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__nand2_2 _3306_ (.A(_2695_),
    .B(_2778_),
    .Y(_2840_));
 sky130_fd_sc_hd__clkbuf_2 _3307_ (.A(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__or2_1 _3308_ (.A(_2839_),
    .B(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__o2111a_1 _3309_ (.A1(_2827_),
    .A2(_2829_),
    .B1(_2833_),
    .C1(_2837_),
    .D1(_2842_),
    .X(_2843_));
 sky130_fd_sc_hd__and4_1 _3310_ (.A(_2794_),
    .B(_2810_),
    .C(_2826_),
    .D(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__inv_2 _3311_ (.A(\BitStream_buffer.BS_buffer[123] ),
    .Y(_2845_));
 sky130_fd_sc_hd__and3_1 _3312_ (.A(\BitStream_buffer.pc[6] ),
    .B(\BitStream_buffer.pc[4] ),
    .C(\BitStream_buffer.pc[5] ),
    .X(_2846_));
 sky130_fd_sc_hd__clkbuf_4 _3313_ (.A(_2846_),
    .X(_2847_));
 sky130_fd_sc_hd__nand2_2 _3314_ (.A(_2620_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__clkbuf_4 _3315_ (.A(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__inv_2 _3316_ (.A(\BitStream_buffer.BS_buffer[121] ),
    .Y(_2850_));
 sky130_fd_sc_hd__nand2_1 _3317_ (.A(net35),
    .B(_2847_),
    .Y(_2851_));
 sky130_fd_sc_hd__clkbuf_2 _3318_ (.A(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__or2_1 _3319_ (.A(_2850_),
    .B(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__inv_2 _3320_ (.A(_2846_),
    .Y(_2854_));
 sky130_fd_sc_hd__nor2_2 _3321_ (.A(_2854_),
    .B(_2615_),
    .Y(_2855_));
 sky130_fd_sc_hd__buf_4 _3322_ (.A(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__nand2_1 _3323_ (.A(_2856_),
    .B(\BitStream_buffer.BS_buffer[122] ),
    .Y(_2857_));
 sky130_fd_sc_hd__nor2_2 _3324_ (.A(_2854_),
    .B(_2634_),
    .Y(_2858_));
 sky130_fd_sc_hd__buf_4 _3325_ (.A(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__nand2_1 _3326_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[120] ),
    .Y(_2860_));
 sky130_fd_sc_hd__o2111a_1 _3327_ (.A1(_2845_),
    .A2(_2849_),
    .B1(_2853_),
    .C1(_2857_),
    .D1(_2860_),
    .X(_2861_));
 sky130_fd_sc_hd__nor2_2 _3328_ (.A(_2854_),
    .B(_2677_),
    .Y(_2862_));
 sky130_fd_sc_hd__buf_2 _3329_ (.A(_2862_),
    .X(_2863_));
 sky130_fd_sc_hd__and2_1 _3330_ (.A(_2680_),
    .B(_2847_),
    .X(_2864_));
 sky130_fd_sc_hd__clkbuf_2 _3331_ (.A(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__buf_2 _3332_ (.A(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__inv_2 _3333_ (.A(\BitStream_buffer.BS_buffer[117] ),
    .Y(_2867_));
 sky130_fd_sc_hd__nand2_2 _3334_ (.A(_2668_),
    .B(_2847_),
    .Y(_2868_));
 sky130_fd_sc_hd__buf_2 _3335_ (.A(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__inv_2 _3336_ (.A(\BitStream_buffer.BS_buffer[116] ),
    .Y(_2870_));
 sky130_fd_sc_hd__nand2_2 _3337_ (.A(_2673_),
    .B(_2847_),
    .Y(_2871_));
 sky130_fd_sc_hd__buf_2 _3338_ (.A(_2871_),
    .X(_2872_));
 sky130_fd_sc_hd__o22ai_1 _3339_ (.A1(_2867_),
    .A2(_2869_),
    .B1(_2870_),
    .B2(_2872_),
    .Y(_2873_));
 sky130_fd_sc_hd__a221oi_1 _3340_ (.A1(\BitStream_buffer.BS_buffer[118] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[119] ),
    .B2(_2866_),
    .C1(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__nor2_2 _3341_ (.A(_2854_),
    .B(_2687_),
    .Y(_2875_));
 sky130_fd_sc_hd__buf_2 _3342_ (.A(_2875_),
    .X(_2876_));
 sky130_fd_sc_hd__and2_1 _3343_ (.A(_2690_),
    .B(_2847_),
    .X(_2877_));
 sky130_fd_sc_hd__clkbuf_2 _3344_ (.A(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__buf_2 _3345_ (.A(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__inv_2 _3346_ (.A(\BitStream_buffer.BS_buffer[125] ),
    .Y(_2880_));
 sky130_fd_sc_hd__nand2_2 _3347_ (.A(_2695_),
    .B(_2847_),
    .Y(_2881_));
 sky130_fd_sc_hd__buf_2 _3348_ (.A(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__inv_2 _3349_ (.A(\BitStream_buffer.BS_buffer[124] ),
    .Y(_2883_));
 sky130_fd_sc_hd__nand2_2 _3350_ (.A(_2700_),
    .B(_2847_),
    .Y(_2884_));
 sky130_fd_sc_hd__buf_2 _3351_ (.A(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__o22ai_1 _3352_ (.A1(_2880_),
    .A2(_2882_),
    .B1(_2883_),
    .B2(_2885_),
    .Y(_2886_));
 sky130_fd_sc_hd__a221oi_1 _3353_ (.A1(\BitStream_buffer.BS_buffer[126] ),
    .A2(_2876_),
    .B1(\BitStream_buffer.BS_buffer[127] ),
    .B2(_2879_),
    .C1(_2886_),
    .Y(_2887_));
 sky130_fd_sc_hd__inv_2 _3354_ (.A(\BitStream_buffer.BS_buffer[112] ),
    .Y(_2888_));
 sky130_fd_sc_hd__nand2_2 _3355_ (.A(_2644_),
    .B(_2847_),
    .Y(_2889_));
 sky130_fd_sc_hd__buf_2 _3356_ (.A(_2889_),
    .X(_2890_));
 sky130_fd_sc_hd__nor2_2 _3357_ (.A(_2854_),
    .B(_2648_),
    .Y(_2891_));
 sky130_fd_sc_hd__buf_2 _3358_ (.A(_2891_),
    .X(_2892_));
 sky130_fd_sc_hd__nand2_1 _3359_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[114] ),
    .Y(_2893_));
 sky130_fd_sc_hd__inv_2 _3360_ (.A(\BitStream_buffer.BS_buffer[115] ),
    .Y(_2894_));
 sky130_fd_sc_hd__nand2_1 _3361_ (.A(_2659_),
    .B(_2846_),
    .Y(_2895_));
 sky130_fd_sc_hd__clkbuf_2 _3362_ (.A(_2895_),
    .X(_2896_));
 sky130_fd_sc_hd__or2_1 _3363_ (.A(_2894_),
    .B(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__inv_2 _3364_ (.A(\BitStream_buffer.BS_buffer[113] ),
    .Y(_2898_));
 sky130_fd_sc_hd__nand2_1 _3365_ (.A(_2654_),
    .B(_2847_),
    .Y(_2899_));
 sky130_fd_sc_hd__clkbuf_2 _3366_ (.A(_2899_),
    .X(_2900_));
 sky130_fd_sc_hd__or2_1 _3367_ (.A(_2898_),
    .B(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__o2111a_1 _3368_ (.A1(_2888_),
    .A2(_2890_),
    .B1(_2893_),
    .C1(_2897_),
    .D1(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__and4_1 _3369_ (.A(_2861_),
    .B(_2874_),
    .C(_2887_),
    .D(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__and4_1 _3370_ (.A(_2705_),
    .B(_2774_),
    .C(_2844_),
    .D(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__inv_2 _3371_ (.A(\BitStream_buffer.BS_buffer[37] ),
    .Y(_2905_));
 sky130_fd_sc_hd__and3_1 _3372_ (.A(_2708_),
    .B(_2600_),
    .C(\BitStream_buffer.pc[5] ),
    .X(_2906_));
 sky130_fd_sc_hd__clkbuf_4 _3373_ (.A(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__nand2_2 _3374_ (.A(_2668_),
    .B(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__clkbuf_4 _3375_ (.A(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__inv_2 _3376_ (.A(\BitStream_buffer.BS_buffer[36] ),
    .Y(_2910_));
 sky130_fd_sc_hd__nand2_2 _3377_ (.A(_2673_),
    .B(_2907_),
    .Y(_2911_));
 sky130_fd_sc_hd__buf_4 _3378_ (.A(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__o22ai_1 _3379_ (.A1(_2905_),
    .A2(_2909_),
    .B1(_2910_),
    .B2(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__inv_2 _3380_ (.A(\BitStream_buffer.BS_buffer[35] ),
    .Y(_2914_));
 sky130_fd_sc_hd__nand2_2 _3381_ (.A(_2659_),
    .B(_2907_),
    .Y(_2915_));
 sky130_fd_sc_hd__buf_2 _3382_ (.A(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__inv_2 _3383_ (.A(\BitStream_buffer.BS_buffer[34] ),
    .Y(_2917_));
 sky130_fd_sc_hd__inv_2 _3384_ (.A(_2648_),
    .Y(_2918_));
 sky130_fd_sc_hd__nand2_2 _3385_ (.A(_2918_),
    .B(_2907_),
    .Y(_2919_));
 sky130_fd_sc_hd__buf_4 _3386_ (.A(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__o22ai_1 _3387_ (.A1(_2914_),
    .A2(_2916_),
    .B1(_2917_),
    .B2(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__inv_2 _3388_ (.A(_2906_),
    .Y(_2922_));
 sky130_fd_sc_hd__nor2_2 _3389_ (.A(_2922_),
    .B(_2677_),
    .Y(_2923_));
 sky130_fd_sc_hd__clkbuf_4 _3390_ (.A(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__and2_2 _3391_ (.A(_2680_),
    .B(_2906_),
    .X(_2925_));
 sky130_fd_sc_hd__clkbuf_4 _3392_ (.A(_2925_),
    .X(_2926_));
 sky130_fd_sc_hd__a22o_1 _3393_ (.A1(\BitStream_buffer.BS_buffer[38] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[39] ),
    .X(_2927_));
 sky130_fd_sc_hd__nor2_2 _3394_ (.A(_2922_),
    .B(_2643_),
    .Y(_2928_));
 sky130_fd_sc_hd__buf_2 _3395_ (.A(_2928_),
    .X(_2929_));
 sky130_fd_sc_hd__and2_2 _3396_ (.A(_2654_),
    .B(_2906_),
    .X(_2930_));
 sky130_fd_sc_hd__clkbuf_4 _3397_ (.A(_2930_),
    .X(_2931_));
 sky130_fd_sc_hd__a22o_1 _3398_ (.A1(\BitStream_buffer.BS_buffer[32] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[33] ),
    .X(_2932_));
 sky130_fd_sc_hd__or4_1 _3399_ (.A(_2913_),
    .B(_2921_),
    .C(_2927_),
    .D(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__nor2_2 _3400_ (.A(_2922_),
    .B(_2699_),
    .Y(_2934_));
 sky130_fd_sc_hd__clkbuf_4 _3401_ (.A(_2934_),
    .X(_2935_));
 sky130_fd_sc_hd__and2_1 _3402_ (.A(_2695_),
    .B(_2907_),
    .X(_2936_));
 sky130_fd_sc_hd__clkbuf_2 _3403_ (.A(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__clkbuf_4 _3404_ (.A(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__inv_2 _3405_ (.A(\BitStream_buffer.BS_buffer[47] ),
    .Y(_2939_));
 sky130_fd_sc_hd__nand2_2 _3406_ (.A(_2690_),
    .B(_2907_),
    .Y(_2940_));
 sky130_fd_sc_hd__buf_2 _3407_ (.A(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__inv_2 _3408_ (.A(\BitStream_buffer.BS_buffer[46] ),
    .Y(_2942_));
 sky130_fd_sc_hd__inv_2 _3409_ (.A(_2687_),
    .Y(_2943_));
 sky130_fd_sc_hd__nand2_2 _3410_ (.A(_2943_),
    .B(_2907_),
    .Y(_2944_));
 sky130_fd_sc_hd__buf_2 _3411_ (.A(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__o22ai_1 _3412_ (.A1(_2939_),
    .A2(_2941_),
    .B1(_2942_),
    .B2(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__a221oi_2 _3413_ (.A1(\BitStream_buffer.BS_buffer[44] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[45] ),
    .B2(_2938_),
    .C1(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__nor2_2 _3414_ (.A(_2922_),
    .B(_2634_),
    .Y(_2948_));
 sky130_fd_sc_hd__buf_2 _3415_ (.A(_2948_),
    .X(_2949_));
 sky130_fd_sc_hd__and2_1 _3416_ (.A(_2628_),
    .B(_2907_),
    .X(_2950_));
 sky130_fd_sc_hd__clkbuf_2 _3417_ (.A(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__buf_2 _3418_ (.A(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__inv_2 _3419_ (.A(\BitStream_buffer.BS_buffer[43] ),
    .Y(_2953_));
 sky130_fd_sc_hd__nand2_2 _3420_ (.A(net36),
    .B(_2907_),
    .Y(_2954_));
 sky130_fd_sc_hd__buf_2 _3421_ (.A(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__inv_2 _3422_ (.A(\BitStream_buffer.BS_buffer[42] ),
    .Y(_2956_));
 sky130_fd_sc_hd__inv_2 _3423_ (.A(_2615_),
    .Y(_2957_));
 sky130_fd_sc_hd__nand2_2 _3424_ (.A(_2957_),
    .B(_2907_),
    .Y(_2958_));
 sky130_fd_sc_hd__clkbuf_4 _3425_ (.A(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__o22ai_1 _3426_ (.A1(_2953_),
    .A2(_2955_),
    .B1(_2956_),
    .B2(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__a221oi_1 _3427_ (.A1(\BitStream_buffer.BS_buffer[40] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[41] ),
    .B2(_2952_),
    .C1(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hd__nand3b_1 _3428_ (.A_N(_2933_),
    .B(_2947_),
    .C(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__inv_2 _3429_ (.A(\BitStream_buffer.BS_buffer[53] ),
    .Y(_2963_));
 sky130_fd_sc_hd__and3_1 _3430_ (.A(_2708_),
    .B(\BitStream_buffer.pc[4] ),
    .C(\BitStream_buffer.pc[5] ),
    .X(_2964_));
 sky130_fd_sc_hd__clkbuf_4 _3431_ (.A(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__nand2_2 _3432_ (.A(_2668_),
    .B(_2965_),
    .Y(_2966_));
 sky130_fd_sc_hd__buf_2 _3433_ (.A(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__inv_2 _3434_ (.A(\BitStream_buffer.BS_buffer[52] ),
    .Y(_2968_));
 sky130_fd_sc_hd__nand2_2 _3435_ (.A(_2673_),
    .B(_2965_),
    .Y(_2969_));
 sky130_fd_sc_hd__buf_4 _3436_ (.A(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__o22ai_1 _3437_ (.A1(_2963_),
    .A2(_2967_),
    .B1(_2968_),
    .B2(_2970_),
    .Y(_2971_));
 sky130_fd_sc_hd__inv_2 _3438_ (.A(\BitStream_buffer.BS_buffer[51] ),
    .Y(_2972_));
 sky130_fd_sc_hd__nand2_2 _3439_ (.A(_2659_),
    .B(_2965_),
    .Y(_2973_));
 sky130_fd_sc_hd__clkbuf_4 _3440_ (.A(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__inv_2 _3441_ (.A(\BitStream_buffer.BS_buffer[50] ),
    .Y(_2975_));
 sky130_fd_sc_hd__nand2_2 _3442_ (.A(_2918_),
    .B(_2965_),
    .Y(_2976_));
 sky130_fd_sc_hd__buf_4 _3443_ (.A(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__o22ai_1 _3444_ (.A1(_2972_),
    .A2(_2974_),
    .B1(_2975_),
    .B2(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__inv_2 _3445_ (.A(_2964_),
    .Y(_2979_));
 sky130_fd_sc_hd__nor2_2 _3446_ (.A(_2979_),
    .B(_2677_),
    .Y(_2980_));
 sky130_fd_sc_hd__clkbuf_4 _3447_ (.A(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__and2_2 _3448_ (.A(_2680_),
    .B(_2964_),
    .X(_2982_));
 sky130_fd_sc_hd__clkbuf_4 _3449_ (.A(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__a22o_1 _3450_ (.A1(\BitStream_buffer.BS_buffer[54] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[55] ),
    .X(_2984_));
 sky130_fd_sc_hd__nor2_2 _3451_ (.A(_2979_),
    .B(_2643_),
    .Y(_2985_));
 sky130_fd_sc_hd__clkbuf_4 _3452_ (.A(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__and2_2 _3453_ (.A(_2654_),
    .B(_2964_),
    .X(_2987_));
 sky130_fd_sc_hd__buf_2 _3454_ (.A(_2987_),
    .X(_2988_));
 sky130_fd_sc_hd__a22o_1 _3455_ (.A1(\BitStream_buffer.BS_buffer[48] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[49] ),
    .X(_2989_));
 sky130_fd_sc_hd__or4_1 _3456_ (.A(_2971_),
    .B(_2978_),
    .C(_2984_),
    .D(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__nor2_2 _3457_ (.A(_2979_),
    .B(_2634_),
    .Y(_2991_));
 sky130_fd_sc_hd__clkbuf_4 _3458_ (.A(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__and2_1 _3459_ (.A(_2628_),
    .B(_2965_),
    .X(_2993_));
 sky130_fd_sc_hd__clkbuf_2 _3460_ (.A(_2993_),
    .X(_2994_));
 sky130_fd_sc_hd__buf_2 _3461_ (.A(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__inv_2 _3462_ (.A(\BitStream_buffer.BS_buffer[59] ),
    .Y(_2996_));
 sky130_fd_sc_hd__nand2_2 _3463_ (.A(net36),
    .B(_2965_),
    .Y(_2997_));
 sky130_fd_sc_hd__buf_2 _3464_ (.A(_2997_),
    .X(_2998_));
 sky130_fd_sc_hd__inv_2 _3465_ (.A(\BitStream_buffer.BS_buffer[58] ),
    .Y(_2999_));
 sky130_fd_sc_hd__nand2_2 _3466_ (.A(_2957_),
    .B(_2965_),
    .Y(_3000_));
 sky130_fd_sc_hd__buf_2 _3467_ (.A(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__o22ai_1 _3468_ (.A1(_2996_),
    .A2(_2998_),
    .B1(_2999_),
    .B2(_3001_),
    .Y(_3002_));
 sky130_fd_sc_hd__a221oi_1 _3469_ (.A1(\BitStream_buffer.BS_buffer[56] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[57] ),
    .B2(_2995_),
    .C1(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__nor2_2 _3470_ (.A(_2979_),
    .B(_2699_),
    .Y(_3004_));
 sky130_fd_sc_hd__buf_2 _3471_ (.A(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__and2_1 _3472_ (.A(_2695_),
    .B(_2965_),
    .X(_3006_));
 sky130_fd_sc_hd__clkbuf_2 _3473_ (.A(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__clkbuf_4 _3474_ (.A(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__inv_2 _3475_ (.A(\BitStream_buffer.BS_buffer[62] ),
    .Y(_3009_));
 sky130_fd_sc_hd__nand2_1 _3476_ (.A(_2943_),
    .B(_2965_),
    .Y(_3010_));
 sky130_fd_sc_hd__clkbuf_2 _3477_ (.A(_3010_),
    .X(_3011_));
 sky130_fd_sc_hd__nand2_2 _3478_ (.A(_2690_),
    .B(_2965_),
    .Y(_3012_));
 sky130_fd_sc_hd__inv_2 _3479_ (.A(_3012_),
    .Y(_3013_));
 sky130_fd_sc_hd__clkbuf_2 _3480_ (.A(_3013_),
    .X(_3014_));
 sky130_fd_sc_hd__a2bb2o_1 _3481_ (.A1_N(_3009_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[63] ),
    .B2(_3014_),
    .X(_3015_));
 sky130_fd_sc_hd__a221oi_1 _3482_ (.A1(\BitStream_buffer.BS_buffer[60] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[61] ),
    .B2(_3008_),
    .C1(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__nand3b_1 _3483_ (.A_N(_2990_),
    .B(_3003_),
    .C(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__inv_2 _3484_ (.A(\BitStream_buffer.BS_buffer[1] ),
    .Y(_3018_));
 sky130_fd_sc_hd__and3_1 _3485_ (.A(_2708_),
    .B(_2600_),
    .C(_2601_),
    .X(_3019_));
 sky130_fd_sc_hd__clkbuf_4 _3486_ (.A(_3019_),
    .X(_3020_));
 sky130_fd_sc_hd__nand2_2 _3487_ (.A(_2654_),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__buf_4 _3488_ (.A(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__nor2_1 _3489_ (.A(_3018_),
    .B(_3022_),
    .Y(_3023_));
 sky130_fd_sc_hd__inv_2 _3490_ (.A(\BitStream_buffer.BS_buffer[7] ),
    .Y(_3024_));
 sky130_fd_sc_hd__nand2_2 _3491_ (.A(_2680_),
    .B(_3020_),
    .Y(_3025_));
 sky130_fd_sc_hd__buf_4 _3492_ (.A(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__inv_2 _3493_ (.A(\BitStream_buffer.BS_buffer[6] ),
    .Y(_3027_));
 sky130_fd_sc_hd__inv_2 _3494_ (.A(_2677_),
    .Y(_3028_));
 sky130_fd_sc_hd__nand2_2 _3495_ (.A(_3028_),
    .B(_3020_),
    .Y(_3029_));
 sky130_fd_sc_hd__buf_4 _3496_ (.A(_3029_),
    .X(_3030_));
 sky130_fd_sc_hd__o22ai_1 _3497_ (.A1(_3024_),
    .A2(_3026_),
    .B1(_3027_),
    .B2(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__inv_2 _3498_ (.A(_3019_),
    .Y(_3032_));
 sky130_fd_sc_hd__nor2_2 _3499_ (.A(_3032_),
    .B(_2672_),
    .Y(_3033_));
 sky130_fd_sc_hd__buf_2 _3500_ (.A(_3033_),
    .X(_3034_));
 sky130_fd_sc_hd__and2_2 _3501_ (.A(_2668_),
    .B(_3020_),
    .X(_3035_));
 sky130_fd_sc_hd__buf_2 _3502_ (.A(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__clkbuf_4 _3503_ (.A(\BitStream_buffer.BS_buffer[5] ),
    .X(_3037_));
 sky130_fd_sc_hd__a22o_1 _3504_ (.A1(\BitStream_buffer.BS_buffer[4] ),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__clkbuf_4 _3505_ (.A(\BitStream_buffer.BS_buffer[2] ),
    .X(_3039_));
 sky130_fd_sc_hd__nor2_2 _3506_ (.A(_3032_),
    .B(_2648_),
    .Y(_3040_));
 sky130_fd_sc_hd__buf_2 _3507_ (.A(_3040_),
    .X(_3041_));
 sky130_fd_sc_hd__and2_2 _3508_ (.A(_2659_),
    .B(_3020_),
    .X(_3042_));
 sky130_fd_sc_hd__clkbuf_4 _3509_ (.A(_3042_),
    .X(_3043_));
 sky130_fd_sc_hd__clkbuf_4 _3510_ (.A(\BitStream_buffer.BS_buffer[3] ),
    .X(_3044_));
 sky130_fd_sc_hd__a22o_1 _3511_ (.A1(_3039_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_3044_),
    .X(_3045_));
 sky130_fd_sc_hd__or4_1 _3512_ (.A(_3023_),
    .B(_3031_),
    .C(_3038_),
    .D(_3045_),
    .X(_3046_));
 sky130_fd_sc_hd__nor2_2 _3513_ (.A(_3032_),
    .B(_2699_),
    .Y(_3047_));
 sky130_fd_sc_hd__buf_2 _3514_ (.A(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__and2_2 _3515_ (.A(_2695_),
    .B(_3019_),
    .X(_3049_));
 sky130_fd_sc_hd__buf_2 _3516_ (.A(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__clkbuf_4 _3517_ (.A(\BitStream_buffer.BS_buffer[13] ),
    .X(_3051_));
 sky130_fd_sc_hd__a22o_1 _3518_ (.A1(\BitStream_buffer.BS_buffer[12] ),
    .A2(_3048_),
    .B1(_3050_),
    .B2(_3051_),
    .X(_3052_));
 sky130_fd_sc_hd__inv_2 _3519_ (.A(\BitStream_buffer.BS_buffer[15] ),
    .Y(_3053_));
 sky130_fd_sc_hd__nand2_2 _3520_ (.A(_2690_),
    .B(_3020_),
    .Y(_3054_));
 sky130_fd_sc_hd__buf_2 _3521_ (.A(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__inv_2 _3522_ (.A(\BitStream_buffer.BS_buffer[14] ),
    .Y(_3056_));
 sky130_fd_sc_hd__nand2_2 _3523_ (.A(_2943_),
    .B(_3020_),
    .Y(_3057_));
 sky130_fd_sc_hd__buf_2 _3524_ (.A(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__o22ai_1 _3525_ (.A1(_3053_),
    .A2(_3055_),
    .B1(_3056_),
    .B2(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__inv_2 _3526_ (.A(\BitStream_buffer.BS_buffer[11] ),
    .Y(_3060_));
 sky130_fd_sc_hd__nand2_2 _3527_ (.A(net36),
    .B(_3020_),
    .Y(_3061_));
 sky130_fd_sc_hd__buf_2 _3528_ (.A(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__inv_2 _3529_ (.A(\BitStream_buffer.BS_buffer[10] ),
    .Y(_3063_));
 sky130_fd_sc_hd__nand2_2 _3530_ (.A(_2957_),
    .B(_3020_),
    .Y(_0322_));
 sky130_fd_sc_hd__buf_2 _3531_ (.A(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__o22ai_1 _3532_ (.A1(_3060_),
    .A2(_3062_),
    .B1(_3063_),
    .B2(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__buf_2 _3533_ (.A(\BitStream_buffer.BS_buffer[9] ),
    .X(_0325_));
 sky130_fd_sc_hd__and2_2 _3534_ (.A(_2628_),
    .B(_3020_),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_4 _3535_ (.A(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_2 _3536_ (.A(_3032_),
    .B(_2634_),
    .Y(_0328_));
 sky130_fd_sc_hd__buf_2 _3537_ (.A(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_4 _3538_ (.A(\BitStream_buffer.BS_buffer[8] ),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _3539_ (.A1(_0325_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__or4_1 _3540_ (.A(_3052_),
    .B(_3059_),
    .C(_0324_),
    .D(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nor2_1 _3541_ (.A(_3046_),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__and3_1 _3542_ (.A(_2708_),
    .B(_2601_),
    .C(\BitStream_buffer.pc[4] ),
    .X(_0334_));
 sky130_fd_sc_hd__inv_2 _3543_ (.A(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nor2_2 _3544_ (.A(_0335_),
    .B(_2634_),
    .Y(_0336_));
 sky130_fd_sc_hd__buf_2 _3545_ (.A(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_4 _3546_ (.A(_0334_),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _3547_ (.A(_2628_),
    .B(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_2 _3548_ (.A(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_4 _3549_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__inv_2 _3550_ (.A(\BitStream_buffer.BS_buffer[27] ),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_2 _3551_ (.A(net36),
    .B(_0338_),
    .Y(_0343_));
 sky130_fd_sc_hd__buf_2 _3552_ (.A(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__inv_2 _3553_ (.A(\BitStream_buffer.BS_buffer[26] ),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_2 _3554_ (.A(_2957_),
    .B(_0338_),
    .Y(_0346_));
 sky130_fd_sc_hd__buf_2 _3555_ (.A(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__o22ai_1 _3556_ (.A1(_0342_),
    .A2(_0344_),
    .B1(_0345_),
    .B2(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__a221oi_1 _3557_ (.A1(\BitStream_buffer.BS_buffer[24] ),
    .A2(_0337_),
    .B1(\BitStream_buffer.BS_buffer[25] ),
    .B2(_0341_),
    .C1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nor2_2 _3558_ (.A(_0335_),
    .B(_2672_),
    .Y(_0350_));
 sky130_fd_sc_hd__buf_2 _3559_ (.A(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__and2_1 _3560_ (.A(_2668_),
    .B(_0338_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_2 _3561_ (.A(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_4 _3562_ (.A(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__inv_2 _3563_ (.A(\BitStream_buffer.BS_buffer[23] ),
    .Y(_0355_));
 sky130_fd_sc_hd__nand2_2 _3564_ (.A(_2680_),
    .B(_0338_),
    .Y(_0356_));
 sky130_fd_sc_hd__buf_2 _3565_ (.A(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__inv_2 _3566_ (.A(\BitStream_buffer.BS_buffer[22] ),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_2 _3567_ (.A(_3028_),
    .B(_0338_),
    .Y(_0359_));
 sky130_fd_sc_hd__buf_2 _3568_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__o22ai_1 _3569_ (.A1(_0355_),
    .A2(_0357_),
    .B1(_0358_),
    .B2(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__a221oi_1 _3570_ (.A1(\BitStream_buffer.BS_buffer[20] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[21] ),
    .B2(_0354_),
    .C1(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__buf_2 _3571_ (.A(\BitStream_buffer.BS_buffer[16] ),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_2 _3572_ (.A(_0335_),
    .B(_2643_),
    .Y(_0364_));
 sky130_fd_sc_hd__buf_2 _3573_ (.A(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_2 _3574_ (.A(\BitStream_buffer.BS_buffer[17] ),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _3575_ (.A(_2654_),
    .B(_0334_),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_2 _3576_ (.A(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__buf_2 _3577_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__inv_2 _3578_ (.A(\BitStream_buffer.BS_buffer[19] ),
    .Y(_0370_));
 sky130_fd_sc_hd__nand2_2 _3579_ (.A(_2659_),
    .B(_0338_),
    .Y(_0371_));
 sky130_fd_sc_hd__buf_2 _3580_ (.A(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__inv_2 _3581_ (.A(\BitStream_buffer.BS_buffer[18] ),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_2 _3582_ (.A(_2918_),
    .B(_0338_),
    .Y(_0374_));
 sky130_fd_sc_hd__buf_2 _3583_ (.A(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__o22ai_1 _3584_ (.A1(_0370_),
    .A2(_0372_),
    .B1(_0373_),
    .B2(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__a221oi_1 _3585_ (.A1(_0363_),
    .A2(_0365_),
    .B1(_0366_),
    .B2(_0369_),
    .C1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_2 _3586_ (.A(_0335_),
    .B(_2699_),
    .Y(_0378_));
 sky130_fd_sc_hd__clkbuf_4 _3587_ (.A(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_4 _3588_ (.A(\BitStream_buffer.BS_buffer[29] ),
    .X(_0380_));
 sky130_fd_sc_hd__and2_1 _3589_ (.A(_2695_),
    .B(_0334_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_2 _3590_ (.A(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_4 _3591_ (.A(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__inv_2 _3592_ (.A(\BitStream_buffer.BS_buffer[31] ),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_2 _3593_ (.A(_2690_),
    .B(_0338_),
    .Y(_0385_));
 sky130_fd_sc_hd__buf_2 _3594_ (.A(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_4 _3595_ (.A(\BitStream_buffer.BS_buffer[30] ),
    .X(_0387_));
 sky130_fd_sc_hd__inv_2 _3596_ (.A(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__nand2_2 _3597_ (.A(_2943_),
    .B(_0338_),
    .Y(_0389_));
 sky130_fd_sc_hd__buf_2 _3598_ (.A(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__o22ai_1 _3599_ (.A1(_0384_),
    .A2(_0386_),
    .B1(_0388_),
    .B2(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__a221oi_1 _3600_ (.A1(\BitStream_buffer.BS_buffer[28] ),
    .A2(_0379_),
    .B1(_0380_),
    .B2(_0383_),
    .C1(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__and4_1 _3601_ (.A(_0349_),
    .B(_0362_),
    .C(_0377_),
    .D(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _3602_ (.A(_0333_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__nor3_1 _3603_ (.A(_2962_),
    .B(_3017_),
    .C(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__a41o_1 _3604_ (.A1(_2612_),
    .A2(_2665_),
    .A3(_2604_),
    .A4(_2626_),
    .B1(_3032_),
    .X(_0396_));
 sky130_fd_sc_hd__and4_1 _3605_ (.A(_0396_),
    .B(_2708_),
    .C(_2600_),
    .D(_2601_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_2 _3606_ (.A(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_2 _3607_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_4 _3608_ (.A(\BitStream_buffer.BS_buffer[0] ),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _3609_ (.A(_0399_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand3_1 _3610_ (.A(_2904_),
    .B(_0395_),
    .C(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _3611_ (.A(\BitStream_buffer.BitStream_buffer_valid_n ),
    .Y(_0403_));
 sky130_fd_sc_hd__buf_4 _3612_ (.A(net19),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_4 _3613_ (.A(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__o21a_1 _3614_ (.A1(\BitStream_buffer.BitStream_buffer_output[15] ),
    .A2(_0403_),
    .B1(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__o21a_1 _3615_ (.A1(_2599_),
    .A2(_0402_),
    .B1(_0406_),
    .X(_0321_));
 sky130_fd_sc_hd__inv_2 _3616_ (.A(\BitStream_buffer.BS_buffer[74] ),
    .Y(_0407_));
 sky130_fd_sc_hd__o22ai_1 _3617_ (.A1(_0407_),
    .A2(_2630_),
    .B1(_2625_),
    .B2(_2637_),
    .Y(_0408_));
 sky130_fd_sc_hd__a221oi_1 _3618_ (.A1(\BitStream_buffer.BS_buffer[75] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[76] ),
    .B2(_2624_),
    .C1(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__nand2_1 _3619_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[67] ),
    .Y(_0410_));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(\BitStream_buffer.BS_buffer[66] ),
    .Y(_0411_));
 sky130_fd_sc_hd__or2_1 _3621_ (.A(_0411_),
    .B(_2656_),
    .X(_0412_));
 sky130_fd_sc_hd__or2_1 _3622_ (.A(_2671_),
    .B(_2661_),
    .X(_0413_));
 sky130_fd_sc_hd__o2111a_1 _3623_ (.A1(_2652_),
    .A2(_2646_),
    .B1(_0410_),
    .C1(_0412_),
    .D1(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__inv_2 _3624_ (.A(\BitStream_buffer.BS_buffer[70] ),
    .Y(_0415_));
 sky130_fd_sc_hd__o22ai_1 _3625_ (.A1(_0415_),
    .A2(_2670_),
    .B1(_2664_),
    .B2(_2675_),
    .Y(_0416_));
 sky130_fd_sc_hd__a22o_1 _3626_ (.A1(\BitStream_buffer.BS_buffer[71] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[72] ),
    .X(_0417_));
 sky130_fd_sc_hd__nor2_1 _3627_ (.A(_0416_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__inv_2 _3628_ (.A(\BitStream_buffer.BS_buffer[78] ),
    .Y(_0419_));
 sky130_fd_sc_hd__o22ai_1 _3629_ (.A1(_0419_),
    .A2(_2697_),
    .B1(_2694_),
    .B2(_2702_),
    .Y(_0420_));
 sky130_fd_sc_hd__a221oi_1 _3630_ (.A1(\BitStream_buffer.BS_buffer[79] ),
    .A2(_2689_),
    .B1(\BitStream_buffer.BS_buffer[80] ),
    .B2(_2693_),
    .C1(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__and4_1 _3631_ (.A(_0409_),
    .B(_0414_),
    .C(_0418_),
    .D(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__inv_2 _3632_ (.A(_2721_),
    .Y(_0423_));
 sky130_fd_sc_hd__or2_1 _3633_ (.A(_2737_),
    .B(_2717_),
    .X(_0424_));
 sky130_fd_sc_hd__nand2_1 _3634_ (.A(_2720_),
    .B(_2714_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand2_1 _3635_ (.A(_2724_),
    .B(_2706_),
    .Y(_0426_));
 sky130_fd_sc_hd__o2111a_1 _3636_ (.A1(_0423_),
    .A2(_2713_),
    .B1(_0424_),
    .C1(_0425_),
    .D1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__inv_2 _3637_ (.A(\BitStream_buffer.BS_buffer[94] ),
    .Y(_0428_));
 sky130_fd_sc_hd__o22ai_1 _3638_ (.A1(_0428_),
    .A2(_2735_),
    .B1(_2733_),
    .B2(_2739_),
    .Y(_0429_));
 sky130_fd_sc_hd__a221oi_1 _3639_ (.A1(\BitStream_buffer.BS_buffer[95] ),
    .A2(_2729_),
    .B1(_2800_),
    .B2(_2732_),
    .C1(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _3640_ (.A(\BitStream_buffer.BS_buffer[82] ),
    .Y(_0431_));
 sky130_fd_sc_hd__nand2_1 _3641_ (.A(_2746_),
    .B(\BitStream_buffer.BS_buffer[83] ),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _3642_ (.A(_2749_),
    .B(\BitStream_buffer.BS_buffer[81] ),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_2 _3643_ (.A(\BitStream_buffer.BS_buffer[84] ),
    .Y(_0434_));
 sky130_fd_sc_hd__or2_1 _3644_ (.A(_0434_),
    .B(_2753_),
    .X(_0435_));
 sky130_fd_sc_hd__o2111a_1 _3645_ (.A1(_0431_),
    .A2(_2744_),
    .B1(_0432_),
    .C1(_0433_),
    .D1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__inv_2 _3646_ (.A(\BitStream_buffer.BS_buffer[88] ),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _3647_ (.A(_2761_),
    .B(_2756_),
    .Y(_0438_));
 sky130_fd_sc_hd__nand2_1 _3648_ (.A(_2765_),
    .B(_2768_),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_2 _3649_ (.A(_2762_),
    .Y(_0440_));
 sky130_fd_sc_hd__or2_1 _3650_ (.A(_0440_),
    .B(_2771_),
    .X(_0441_));
 sky130_fd_sc_hd__o2111a_1 _3651_ (.A1(_0437_),
    .A2(_2759_),
    .B1(_0438_),
    .C1(_0439_),
    .D1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__and4_1 _3652_ (.A(_0427_),
    .B(_0430_),
    .C(_0436_),
    .D(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__inv_2 _3653_ (.A(_2788_),
    .Y(_0444_));
 sky130_fd_sc_hd__inv_2 _3654_ (.A(\BitStream_buffer.BS_buffer[108] ),
    .Y(_0445_));
 sky130_fd_sc_hd__or2_1 _3655_ (.A(_0445_),
    .B(_2784_),
    .X(_0446_));
 sky130_fd_sc_hd__nand2_1 _3656_ (.A(_2787_),
    .B(_2781_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_1 _3657_ (.A(_2791_),
    .B(\BitStream_buffer.BS_buffer[105] ),
    .Y(_0448_));
 sky130_fd_sc_hd__o2111a_1 _3658_ (.A1(_0444_),
    .A2(_2780_),
    .B1(_0446_),
    .C1(_0447_),
    .D1(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__inv_2 _3659_ (.A(_2820_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_1 _3660_ (.A(_2799_),
    .B(\BitStream_buffer.BS_buffer[97] ),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _3661_ (.A(_2803_),
    .B(\BitStream_buffer.BS_buffer[99] ),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _3662_ (.A(_2804_),
    .Y(_0453_));
 sky130_fd_sc_hd__or2_1 _3663_ (.A(_0453_),
    .B(_2808_),
    .X(_0454_));
 sky130_fd_sc_hd__o2111a_1 _3664_ (.A1(_0450_),
    .A2(_2797_),
    .B1(_0451_),
    .C1(_0452_),
    .D1(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__inv_2 _3665_ (.A(_2792_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _3666_ (.A(_2815_),
    .B(\BitStream_buffer.BS_buffer[103] ),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _3667_ (.A(_2819_),
    .B(\BitStream_buffer.BS_buffer[101] ),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _3668_ (.A(_2816_),
    .Y(_0459_));
 sky130_fd_sc_hd__or2_1 _3669_ (.A(_0459_),
    .B(_2824_),
    .X(_0460_));
 sky130_fd_sc_hd__o2111a_1 _3670_ (.A1(_0456_),
    .A2(_2813_),
    .B1(_0457_),
    .C1(_0458_),
    .D1(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _3671_ (.A(_2831_),
    .B(_2838_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _3672_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[111] ),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_2 _3673_ (.A(_2836_),
    .Y(_0464_));
 sky130_fd_sc_hd__or2_1 _3674_ (.A(_0464_),
    .B(_2841_),
    .X(_0465_));
 sky130_fd_sc_hd__o2111a_1 _3675_ (.A1(_2888_),
    .A2(_2829_),
    .B1(_0462_),
    .C1(_0463_),
    .D1(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__and4_1 _3676_ (.A(_0449_),
    .B(_0455_),
    .C(_0461_),
    .D(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__inv_2 _3677_ (.A(\BitStream_buffer.BS_buffer[122] ),
    .Y(_0468_));
 sky130_fd_sc_hd__or2_1 _3678_ (.A(_0468_),
    .B(_2852_),
    .X(_0469_));
 sky130_fd_sc_hd__nand2_1 _3679_ (.A(_2856_),
    .B(\BitStream_buffer.BS_buffer[123] ),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _3680_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[121] ),
    .Y(_0471_));
 sky130_fd_sc_hd__o2111a_1 _3681_ (.A1(_2883_),
    .A2(_2849_),
    .B1(_0469_),
    .C1(_0470_),
    .D1(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__inv_2 _3682_ (.A(\BitStream_buffer.BS_buffer[118] ),
    .Y(_0473_));
 sky130_fd_sc_hd__o22ai_1 _3683_ (.A1(_0473_),
    .A2(_2869_),
    .B1(_2867_),
    .B2(_2872_),
    .Y(_0474_));
 sky130_fd_sc_hd__a221oi_1 _3684_ (.A1(\BitStream_buffer.BS_buffer[119] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[120] ),
    .B2(_2866_),
    .C1(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__inv_2 _3685_ (.A(\BitStream_buffer.BS_buffer[126] ),
    .Y(_0476_));
 sky130_fd_sc_hd__o22ai_1 _3686_ (.A1(_0476_),
    .A2(_2882_),
    .B1(_2880_),
    .B2(_2885_),
    .Y(_0477_));
 sky130_fd_sc_hd__a221oi_1 _3687_ (.A1(_0400_),
    .A2(_2878_),
    .B1(\BitStream_buffer.BS_buffer[127] ),
    .B2(_2876_),
    .C1(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[115] ),
    .Y(_0479_));
 sky130_fd_sc_hd__or2_1 _3689_ (.A(_2870_),
    .B(_2896_),
    .X(_0480_));
 sky130_fd_sc_hd__inv_2 _3690_ (.A(\BitStream_buffer.BS_buffer[114] ),
    .Y(_0481_));
 sky130_fd_sc_hd__or2_1 _3691_ (.A(_0481_),
    .B(_2900_),
    .X(_0482_));
 sky130_fd_sc_hd__o2111a_1 _3692_ (.A1(_2898_),
    .A2(_2890_),
    .B1(_0479_),
    .C1(_0480_),
    .D1(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__and4_1 _3693_ (.A(_0472_),
    .B(_0475_),
    .C(_0478_),
    .D(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__and4_1 _3694_ (.A(_0422_),
    .B(_0443_),
    .C(_0467_),
    .D(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__inv_2 _3695_ (.A(\BitStream_buffer.BS_buffer[38] ),
    .Y(_0486_));
 sky130_fd_sc_hd__o22ai_1 _3696_ (.A1(_0486_),
    .A2(_2909_),
    .B1(_2905_),
    .B2(_2912_),
    .Y(_0487_));
 sky130_fd_sc_hd__o22ai_1 _3697_ (.A1(_2910_),
    .A2(_2916_),
    .B1(_2914_),
    .B2(_2920_),
    .Y(_0488_));
 sky130_fd_sc_hd__a22o_1 _3698_ (.A1(\BitStream_buffer.BS_buffer[39] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[40] ),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _3699_ (.A1(\BitStream_buffer.BS_buffer[33] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[34] ),
    .X(_0490_));
 sky130_fd_sc_hd__or4_1 _3700_ (.A(_0487_),
    .B(_0488_),
    .C(_0489_),
    .D(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__inv_2 _3701_ (.A(\BitStream_buffer.BS_buffer[48] ),
    .Y(_0492_));
 sky130_fd_sc_hd__o22ai_1 _3702_ (.A1(_0492_),
    .A2(_2941_),
    .B1(_2939_),
    .B2(_2945_),
    .Y(_0493_));
 sky130_fd_sc_hd__a221oi_1 _3703_ (.A1(\BitStream_buffer.BS_buffer[45] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[46] ),
    .B2(_2938_),
    .C1(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _3704_ (.A(\BitStream_buffer.BS_buffer[44] ),
    .Y(_0495_));
 sky130_fd_sc_hd__o22ai_1 _3705_ (.A1(_0495_),
    .A2(_2955_),
    .B1(_2953_),
    .B2(_2959_),
    .Y(_0496_));
 sky130_fd_sc_hd__a221oi_1 _3706_ (.A1(\BitStream_buffer.BS_buffer[41] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[42] ),
    .B2(_2952_),
    .C1(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand3b_1 _3707_ (.A_N(_0491_),
    .B(_0494_),
    .C(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _3708_ (.A(\BitStream_buffer.BS_buffer[54] ),
    .Y(_0499_));
 sky130_fd_sc_hd__o22ai_1 _3709_ (.A1(_0499_),
    .A2(_2967_),
    .B1(_2963_),
    .B2(_2970_),
    .Y(_0500_));
 sky130_fd_sc_hd__o22ai_1 _3710_ (.A1(_2968_),
    .A2(_2974_),
    .B1(_2972_),
    .B2(_2977_),
    .Y(_0501_));
 sky130_fd_sc_hd__a22o_1 _3711_ (.A1(\BitStream_buffer.BS_buffer[55] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[56] ),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _3712_ (.A1(\BitStream_buffer.BS_buffer[49] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[50] ),
    .X(_0503_));
 sky130_fd_sc_hd__or4_1 _3713_ (.A(_0500_),
    .B(_0501_),
    .C(_0502_),
    .D(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__inv_2 _3714_ (.A(\BitStream_buffer.BS_buffer[60] ),
    .Y(_0505_));
 sky130_fd_sc_hd__o22ai_1 _3715_ (.A1(_0505_),
    .A2(_2998_),
    .B1(_2996_),
    .B2(_3001_),
    .Y(_0506_));
 sky130_fd_sc_hd__a221oi_1 _3716_ (.A1(\BitStream_buffer.BS_buffer[57] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[58] ),
    .B2(_2995_),
    .C1(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_2 _3717_ (.A(\BitStream_buffer.BS_buffer[63] ),
    .Y(_0508_));
 sky130_fd_sc_hd__a2bb2o_1 _3718_ (.A1_N(_0508_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[64] ),
    .B2(_3014_),
    .X(_0509_));
 sky130_fd_sc_hd__a221oi_1 _3719_ (.A1(\BitStream_buffer.BS_buffer[61] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[62] ),
    .B2(_3008_),
    .C1(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand3b_1 _3720_ (.A_N(_0504_),
    .B(_0507_),
    .C(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _3721_ (.A(_3039_),
    .Y(_0512_));
 sky130_fd_sc_hd__nor2_1 _3722_ (.A(_0512_),
    .B(_3022_),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _3723_ (.A(\BitStream_buffer.BS_buffer[8] ),
    .Y(_0514_));
 sky130_fd_sc_hd__o22ai_1 _3724_ (.A1(_0514_),
    .A2(_3026_),
    .B1(_3024_),
    .B2(_3030_),
    .Y(_0515_));
 sky130_fd_sc_hd__clkbuf_4 _3725_ (.A(\BitStream_buffer.BS_buffer[6] ),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _3726_ (.A1(\BitStream_buffer.BS_buffer[5] ),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_4 _3727_ (.A(\BitStream_buffer.BS_buffer[4] ),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _3728_ (.A1(_3044_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__or4_1 _3729_ (.A(_0513_),
    .B(_0515_),
    .C(_0517_),
    .D(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_4 _3730_ (.A(\BitStream_buffer.BS_buffer[14] ),
    .X(_0521_));
 sky130_fd_sc_hd__a22o_1 _3731_ (.A1(\BitStream_buffer.BS_buffer[13] ),
    .A2(_3048_),
    .B1(_3050_),
    .B2(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__inv_2 _3732_ (.A(\BitStream_buffer.BS_buffer[16] ),
    .Y(_0523_));
 sky130_fd_sc_hd__o22ai_1 _3733_ (.A1(_0523_),
    .A2(_3055_),
    .B1(_3053_),
    .B2(_3058_),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _3734_ (.A(\BitStream_buffer.BS_buffer[12] ),
    .Y(_0525_));
 sky130_fd_sc_hd__o22ai_1 _3735_ (.A1(_0525_),
    .A2(_3062_),
    .B1(_3060_),
    .B2(_0323_),
    .Y(_0526_));
 sky130_fd_sc_hd__clkbuf_4 _3736_ (.A(\BitStream_buffer.BS_buffer[10] ),
    .X(_0527_));
 sky130_fd_sc_hd__a22o_1 _3737_ (.A1(_0527_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0325_),
    .X(_0528_));
 sky130_fd_sc_hd__or4_1 _3738_ (.A(_0522_),
    .B(_0524_),
    .C(_0526_),
    .D(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__nor2_1 _3739_ (.A(_0520_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _3740_ (.A(\BitStream_buffer.BS_buffer[28] ),
    .Y(_0531_));
 sky130_fd_sc_hd__o22ai_1 _3741_ (.A1(_0531_),
    .A2(_0344_),
    .B1(_0342_),
    .B2(_0347_),
    .Y(_0532_));
 sky130_fd_sc_hd__a221oi_1 _3742_ (.A1(\BitStream_buffer.BS_buffer[25] ),
    .A2(_0337_),
    .B1(\BitStream_buffer.BS_buffer[26] ),
    .B2(_0341_),
    .C1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _3743_ (.A(\BitStream_buffer.BS_buffer[24] ),
    .Y(_0534_));
 sky130_fd_sc_hd__o22ai_1 _3744_ (.A1(_0534_),
    .A2(_0357_),
    .B1(_0355_),
    .B2(_0360_),
    .Y(_0535_));
 sky130_fd_sc_hd__a221oi_1 _3745_ (.A1(\BitStream_buffer.BS_buffer[21] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[22] ),
    .B2(_0354_),
    .C1(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_2 _3746_ (.A(\BitStream_buffer.BS_buffer[20] ),
    .Y(_0537_));
 sky130_fd_sc_hd__o22ai_1 _3747_ (.A1(_0537_),
    .A2(_0372_),
    .B1(_0370_),
    .B2(_0375_),
    .Y(_0538_));
 sky130_fd_sc_hd__a221oi_1 _3748_ (.A1(_0366_),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[18] ),
    .B2(_0369_),
    .C1(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__inv_2 _3749_ (.A(\BitStream_buffer.BS_buffer[32] ),
    .Y(_0540_));
 sky130_fd_sc_hd__o22ai_1 _3750_ (.A1(_0540_),
    .A2(_0386_),
    .B1(_0384_),
    .B2(_0390_),
    .Y(_0541_));
 sky130_fd_sc_hd__a221oi_1 _3751_ (.A1(_0380_),
    .A2(_0379_),
    .B1(_0387_),
    .B2(_0383_),
    .C1(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__and4_1 _3752_ (.A(_0533_),
    .B(_0536_),
    .C(_0539_),
    .D(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _3753_ (.A(_0530_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__nor3_1 _3754_ (.A(_0498_),
    .B(_0511_),
    .C(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _3755_ (.A(_0399_),
    .B(\BitStream_buffer.BS_buffer[1] ),
    .Y(_0546_));
 sky130_fd_sc_hd__nand3_1 _3756_ (.A(_0485_),
    .B(_0545_),
    .C(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__o21a_1 _3757_ (.A1(\BitStream_buffer.BitStream_buffer_output[14] ),
    .A2(_0403_),
    .B1(_0405_),
    .X(_0548_));
 sky130_fd_sc_hd__o21a_1 _3758_ (.A1(_2599_),
    .A2(_0547_),
    .B1(_0548_),
    .X(_0320_));
 sky130_fd_sc_hd__inv_2 _3759_ (.A(\BitStream_buffer.BS_buffer[75] ),
    .Y(_0549_));
 sky130_fd_sc_hd__o22ai_1 _3760_ (.A1(_0549_),
    .A2(_2630_),
    .B1(_0407_),
    .B2(_2637_),
    .Y(_0550_));
 sky130_fd_sc_hd__a221oi_1 _3761_ (.A1(\BitStream_buffer.BS_buffer[76] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[77] ),
    .B2(_2624_),
    .C1(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _3762_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[68] ),
    .Y(_0552_));
 sky130_fd_sc_hd__or2_1 _3763_ (.A(_2658_),
    .B(_2656_),
    .X(_0553_));
 sky130_fd_sc_hd__or2_1 _3764_ (.A(_2664_),
    .B(_2661_),
    .X(_0554_));
 sky130_fd_sc_hd__o2111a_1 _3765_ (.A1(_0411_),
    .A2(_2646_),
    .B1(_0552_),
    .C1(_0553_),
    .D1(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__inv_2 _3766_ (.A(\BitStream_buffer.BS_buffer[71] ),
    .Y(_0556_));
 sky130_fd_sc_hd__o22ai_1 _3767_ (.A1(_0556_),
    .A2(_2670_),
    .B1(_0415_),
    .B2(_2675_),
    .Y(_0557_));
 sky130_fd_sc_hd__a22o_1 _3768_ (.A1(\BitStream_buffer.BS_buffer[72] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[73] ),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_1 _3769_ (.A(_0557_),
    .B(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_2 _3770_ (.A(\BitStream_buffer.BS_buffer[79] ),
    .Y(_0560_));
 sky130_fd_sc_hd__o22ai_1 _3771_ (.A1(_0560_),
    .A2(_2697_),
    .B1(_0419_),
    .B2(_2702_),
    .Y(_0561_));
 sky130_fd_sc_hd__a221oi_1 _3772_ (.A1(\BitStream_buffer.BS_buffer[80] ),
    .A2(_2689_),
    .B1(\BitStream_buffer.BS_buffer[81] ),
    .B2(_2693_),
    .C1(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__and4_1 _3773_ (.A(_0551_),
    .B(_0555_),
    .C(_0559_),
    .D(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(_2733_),
    .B(_2717_),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _3775_ (.A(_2720_),
    .B(_2736_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_1 _3776_ (.A(_2724_),
    .B(_2721_),
    .Y(_0566_));
 sky130_fd_sc_hd__o2111a_1 _3777_ (.A1(_2715_),
    .A2(_2713_),
    .B1(_0564_),
    .C1(_0565_),
    .D1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__inv_2 _3778_ (.A(\BitStream_buffer.BS_buffer[95] ),
    .Y(_0568_));
 sky130_fd_sc_hd__o22ai_1 _3779_ (.A1(_0568_),
    .A2(_2735_),
    .B1(_0428_),
    .B2(_2739_),
    .Y(_0569_));
 sky130_fd_sc_hd__a221oi_1 _3780_ (.A1(_2800_),
    .A2(_2729_),
    .B1(\BitStream_buffer.BS_buffer[97] ),
    .B2(_2732_),
    .C1(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_1 _3781_ (.A(_2746_),
    .B(_2766_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_1 _3782_ (.A(_2749_),
    .B(\BitStream_buffer.BS_buffer[82] ),
    .Y(_0572_));
 sky130_fd_sc_hd__or2_1 _3783_ (.A(_2769_),
    .B(_2753_),
    .X(_0573_));
 sky130_fd_sc_hd__o2111a_1 _3784_ (.A1(_2751_),
    .A2(_2744_),
    .B1(_0571_),
    .C1(_0572_),
    .D1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__nand2_1 _3785_ (.A(_2761_),
    .B(_2725_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _3786_ (.A(_2765_),
    .B(_2762_),
    .Y(_0576_));
 sky130_fd_sc_hd__or2_1 _3787_ (.A(_2757_),
    .B(_2771_),
    .X(_0577_));
 sky130_fd_sc_hd__o2111a_1 _3788_ (.A1(_2707_),
    .A2(_2759_),
    .B1(_0575_),
    .C1(_0576_),
    .D1(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__and4_1 _3789_ (.A(_0567_),
    .B(_0570_),
    .C(_0574_),
    .D(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__or2_1 _3790_ (.A(_2839_),
    .B(_2784_),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_1 _3791_ (.A(_2787_),
    .B(_2832_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _3792_ (.A(_2791_),
    .B(_2788_),
    .Y(_0582_));
 sky130_fd_sc_hd__o2111a_1 _3793_ (.A1(_2782_),
    .A2(_2780_),
    .B1(_0580_),
    .C1(_0581_),
    .D1(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _3794_ (.A(_2799_),
    .B(_2804_),
    .Y(_0584_));
 sky130_fd_sc_hd__nand2_1 _3795_ (.A(_2803_),
    .B(_2820_),
    .Y(_0585_));
 sky130_fd_sc_hd__or2_1 _3796_ (.A(_2795_),
    .B(_2808_),
    .X(_0586_));
 sky130_fd_sc_hd__o2111a_1 _3797_ (.A1(_2822_),
    .A2(_2797_),
    .B1(_0584_),
    .C1(_0585_),
    .D1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__nand2_1 _3798_ (.A(_2815_),
    .B(_2792_),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(_2819_),
    .B(_2816_),
    .Y(_0589_));
 sky130_fd_sc_hd__or2_1 _3800_ (.A(_2811_),
    .B(_2824_),
    .X(_0590_));
 sky130_fd_sc_hd__o2111a_1 _3801_ (.A1(_2775_),
    .A2(_2813_),
    .B1(_0588_),
    .C1(_0589_),
    .D1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__nand2_1 _3802_ (.A(_2831_),
    .B(_2836_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _3803_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[112] ),
    .Y(_0593_));
 sky130_fd_sc_hd__or2_1 _3804_ (.A(_2827_),
    .B(_2841_),
    .X(_0594_));
 sky130_fd_sc_hd__o2111a_1 _3805_ (.A1(_2898_),
    .A2(_2829_),
    .B1(_0592_),
    .C1(_0593_),
    .D1(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__and4_1 _3806_ (.A(_0583_),
    .B(_0587_),
    .C(_0591_),
    .D(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__or2_1 _3807_ (.A(_2845_),
    .B(_2852_),
    .X(_0597_));
 sky130_fd_sc_hd__nand2_1 _3808_ (.A(_2856_),
    .B(\BitStream_buffer.BS_buffer[124] ),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2_1 _3809_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[122] ),
    .Y(_0599_));
 sky130_fd_sc_hd__o2111a_1 _3810_ (.A1(_2880_),
    .A2(_2849_),
    .B1(_0597_),
    .C1(_0598_),
    .D1(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__inv_2 _3811_ (.A(\BitStream_buffer.BS_buffer[119] ),
    .Y(_0601_));
 sky130_fd_sc_hd__o22ai_1 _3812_ (.A1(_0601_),
    .A2(_2869_),
    .B1(_0473_),
    .B2(_2872_),
    .Y(_0602_));
 sky130_fd_sc_hd__a221oi_1 _3813_ (.A1(\BitStream_buffer.BS_buffer[120] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[121] ),
    .B2(_2866_),
    .C1(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _3814_ (.A(\BitStream_buffer.BS_buffer[127] ),
    .Y(_0604_));
 sky130_fd_sc_hd__o22ai_1 _3815_ (.A1(_0604_),
    .A2(_2882_),
    .B1(_0476_),
    .B2(_2885_),
    .Y(_0605_));
 sky130_fd_sc_hd__a221oi_1 _3816_ (.A1(_0400_),
    .A2(_2876_),
    .B1(\BitStream_buffer.BS_buffer[1] ),
    .B2(_2879_),
    .C1(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _3817_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[116] ),
    .Y(_0607_));
 sky130_fd_sc_hd__or2_1 _3818_ (.A(_2867_),
    .B(_2896_),
    .X(_0608_));
 sky130_fd_sc_hd__or2_1 _3819_ (.A(_2894_),
    .B(_2900_),
    .X(_0609_));
 sky130_fd_sc_hd__o2111a_1 _3820_ (.A1(_0481_),
    .A2(_2890_),
    .B1(_0607_),
    .C1(_0608_),
    .D1(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__and4_1 _3821_ (.A(_0600_),
    .B(_0603_),
    .C(_0606_),
    .D(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__and4_1 _3822_ (.A(_0563_),
    .B(_0579_),
    .C(_0596_),
    .D(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__inv_2 _3823_ (.A(\BitStream_buffer.BS_buffer[39] ),
    .Y(_0613_));
 sky130_fd_sc_hd__o22ai_1 _3824_ (.A1(_0613_),
    .A2(_2909_),
    .B1(_0486_),
    .B2(_2912_),
    .Y(_0614_));
 sky130_fd_sc_hd__o22ai_1 _3825_ (.A1(_2905_),
    .A2(_2916_),
    .B1(_2910_),
    .B2(_2920_),
    .Y(_0615_));
 sky130_fd_sc_hd__a22o_1 _3826_ (.A1(\BitStream_buffer.BS_buffer[40] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[41] ),
    .X(_0616_));
 sky130_fd_sc_hd__a22o_1 _3827_ (.A1(\BitStream_buffer.BS_buffer[34] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[35] ),
    .X(_0617_));
 sky130_fd_sc_hd__or4_1 _3828_ (.A(_0614_),
    .B(_0615_),
    .C(_0616_),
    .D(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__inv_2 _3829_ (.A(\BitStream_buffer.BS_buffer[49] ),
    .Y(_0619_));
 sky130_fd_sc_hd__o22ai_1 _3830_ (.A1(_0619_),
    .A2(_2941_),
    .B1(_0492_),
    .B2(_2945_),
    .Y(_0620_));
 sky130_fd_sc_hd__a221oi_1 _3831_ (.A1(\BitStream_buffer.BS_buffer[46] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[47] ),
    .B2(_2938_),
    .C1(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__inv_2 _3832_ (.A(\BitStream_buffer.BS_buffer[45] ),
    .Y(_0622_));
 sky130_fd_sc_hd__o22ai_1 _3833_ (.A1(_0622_),
    .A2(_2955_),
    .B1(_0495_),
    .B2(_2959_),
    .Y(_0623_));
 sky130_fd_sc_hd__a221oi_1 _3834_ (.A1(\BitStream_buffer.BS_buffer[42] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[43] ),
    .B2(_2952_),
    .C1(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand3b_1 _3835_ (.A_N(_0618_),
    .B(_0621_),
    .C(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_2 _3836_ (.A(\BitStream_buffer.BS_buffer[55] ),
    .Y(_0626_));
 sky130_fd_sc_hd__o22ai_1 _3837_ (.A1(_0626_),
    .A2(_2967_),
    .B1(_0499_),
    .B2(_2970_),
    .Y(_0627_));
 sky130_fd_sc_hd__o22ai_1 _3838_ (.A1(_2963_),
    .A2(_2974_),
    .B1(_2968_),
    .B2(_2977_),
    .Y(_0628_));
 sky130_fd_sc_hd__a22o_1 _3839_ (.A1(\BitStream_buffer.BS_buffer[56] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[57] ),
    .X(_0629_));
 sky130_fd_sc_hd__a22o_1 _3840_ (.A1(\BitStream_buffer.BS_buffer[50] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[51] ),
    .X(_0630_));
 sky130_fd_sc_hd__or4_1 _3841_ (.A(_0627_),
    .B(_0628_),
    .C(_0629_),
    .D(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__inv_2 _3842_ (.A(\BitStream_buffer.BS_buffer[61] ),
    .Y(_0632_));
 sky130_fd_sc_hd__o22ai_1 _3843_ (.A1(_0632_),
    .A2(_2998_),
    .B1(_0505_),
    .B2(_3001_),
    .Y(_0633_));
 sky130_fd_sc_hd__a221oi_1 _3844_ (.A1(\BitStream_buffer.BS_buffer[58] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[59] ),
    .B2(_2995_),
    .C1(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__a2bb2o_1 _3845_ (.A1_N(_2640_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[65] ),
    .B2(_3014_),
    .X(_0635_));
 sky130_fd_sc_hd__a221oi_1 _3846_ (.A1(\BitStream_buffer.BS_buffer[62] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[63] ),
    .B2(_3008_),
    .C1(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand3b_1 _3847_ (.A_N(_0631_),
    .B(_0634_),
    .C(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__inv_2 _3848_ (.A(\BitStream_buffer.BS_buffer[3] ),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_1 _3849_ (.A(_0638_),
    .B(_3022_),
    .Y(_0639_));
 sky130_fd_sc_hd__inv_2 _3850_ (.A(\BitStream_buffer.BS_buffer[9] ),
    .Y(_0640_));
 sky130_fd_sc_hd__o22ai_1 _3851_ (.A1(_0640_),
    .A2(_3026_),
    .B1(_0514_),
    .B2(_3030_),
    .Y(_0641_));
 sky130_fd_sc_hd__a22o_1 _3852_ (.A1(_0516_),
    .A2(_3034_),
    .B1(_3036_),
    .B2(\BitStream_buffer.BS_buffer[7] ),
    .X(_0642_));
 sky130_fd_sc_hd__a22o_1 _3853_ (.A1(_0518_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_3037_),
    .X(_0643_));
 sky130_fd_sc_hd__or4_1 _3854_ (.A(_0639_),
    .B(_0641_),
    .C(_0642_),
    .D(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__a22o_1 _3855_ (.A1(_0521_),
    .A2(_3048_),
    .B1(_3050_),
    .B2(\BitStream_buffer.BS_buffer[15] ),
    .X(_0645_));
 sky130_fd_sc_hd__inv_2 _3856_ (.A(\BitStream_buffer.BS_buffer[17] ),
    .Y(_0646_));
 sky130_fd_sc_hd__o22ai_1 _3857_ (.A1(_0646_),
    .A2(_3055_),
    .B1(_0523_),
    .B2(_3058_),
    .Y(_0647_));
 sky130_fd_sc_hd__inv_2 _3858_ (.A(\BitStream_buffer.BS_buffer[13] ),
    .Y(_0648_));
 sky130_fd_sc_hd__o22ai_1 _3859_ (.A1(_0648_),
    .A2(_3062_),
    .B1(_0525_),
    .B2(_0323_),
    .Y(_0649_));
 sky130_fd_sc_hd__clkbuf_4 _3860_ (.A(\BitStream_buffer.BS_buffer[11] ),
    .X(_0650_));
 sky130_fd_sc_hd__a22o_1 _3861_ (.A1(_0650_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0527_),
    .X(_0651_));
 sky130_fd_sc_hd__or4_1 _3862_ (.A(_0645_),
    .B(_0647_),
    .C(_0649_),
    .D(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__nor2_1 _3863_ (.A(_0644_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__inv_2 _3864_ (.A(_0380_),
    .Y(_0654_));
 sky130_fd_sc_hd__o22ai_1 _3865_ (.A1(_0654_),
    .A2(_0344_),
    .B1(_0531_),
    .B2(_0347_),
    .Y(_0655_));
 sky130_fd_sc_hd__a221oi_1 _3866_ (.A1(\BitStream_buffer.BS_buffer[26] ),
    .A2(_0337_),
    .B1(\BitStream_buffer.BS_buffer[27] ),
    .B2(_0341_),
    .C1(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__inv_2 _3867_ (.A(\BitStream_buffer.BS_buffer[25] ),
    .Y(_0657_));
 sky130_fd_sc_hd__o22ai_1 _3868_ (.A1(_0657_),
    .A2(_0357_),
    .B1(_0534_),
    .B2(_0360_),
    .Y(_0658_));
 sky130_fd_sc_hd__a221oi_1 _3869_ (.A1(\BitStream_buffer.BS_buffer[22] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[23] ),
    .B2(_0354_),
    .C1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__inv_2 _3870_ (.A(\BitStream_buffer.BS_buffer[21] ),
    .Y(_0660_));
 sky130_fd_sc_hd__o22ai_1 _3871_ (.A1(_0660_),
    .A2(_0372_),
    .B1(_0537_),
    .B2(_0375_),
    .Y(_0661_));
 sky130_fd_sc_hd__a221oi_1 _3872_ (.A1(\BitStream_buffer.BS_buffer[18] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[19] ),
    .B2(_0369_),
    .C1(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__inv_2 _3873_ (.A(\BitStream_buffer.BS_buffer[33] ),
    .Y(_0663_));
 sky130_fd_sc_hd__o22ai_1 _3874_ (.A1(_0663_),
    .A2(_0386_),
    .B1(_0540_),
    .B2(_0390_),
    .Y(_0664_));
 sky130_fd_sc_hd__a221oi_1 _3875_ (.A1(_0387_),
    .A2(_0379_),
    .B1(\BitStream_buffer.BS_buffer[31] ),
    .B2(_0383_),
    .C1(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__and4_1 _3876_ (.A(_0656_),
    .B(_0659_),
    .C(_0662_),
    .D(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(_0653_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__nor3_1 _3878_ (.A(_0625_),
    .B(_0637_),
    .C(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_1 _3879_ (.A(_0399_),
    .B(_3039_),
    .Y(_0669_));
 sky130_fd_sc_hd__nand3_1 _3880_ (.A(_0612_),
    .B(_0668_),
    .C(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__inv_2 _3881_ (.A(\BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_0671_));
 sky130_fd_sc_hd__buf_2 _3882_ (.A(_2598_),
    .X(_0672_));
 sky130_fd_sc_hd__inv_2 _3883_ (.A(net19),
    .Y(_0673_));
 sky130_fd_sc_hd__buf_2 _3884_ (.A(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_4 _3885_ (.A(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__a21oi_1 _3886_ (.A1(_0671_),
    .A2(_0672_),
    .B1(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__o21a_1 _3887_ (.A1(_2599_),
    .A2(_0670_),
    .B1(_0676_),
    .X(_0319_));
 sky130_fd_sc_hd__o22ai_1 _3888_ (.A1(_2698_),
    .A2(_2630_),
    .B1(_0549_),
    .B2(_2637_),
    .Y(_0677_));
 sky130_fd_sc_hd__a221oi_1 _3889_ (.A1(\BitStream_buffer.BS_buffer[77] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[78] ),
    .B2(_2624_),
    .C1(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _3890_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[69] ),
    .Y(_0679_));
 sky130_fd_sc_hd__or2_1 _3891_ (.A(_2671_),
    .B(_2656_),
    .X(_0680_));
 sky130_fd_sc_hd__or2_1 _3892_ (.A(_0415_),
    .B(_2661_),
    .X(_0681_));
 sky130_fd_sc_hd__o2111a_1 _3893_ (.A1(_2658_),
    .A2(_2646_),
    .B1(_0679_),
    .C1(_0680_),
    .D1(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__o22ai_1 _3894_ (.A1(_2631_),
    .A2(_2670_),
    .B1(_0556_),
    .B2(_2675_),
    .Y(_0683_));
 sky130_fd_sc_hd__a22o_1 _3895_ (.A1(\BitStream_buffer.BS_buffer[73] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[74] ),
    .X(_0684_));
 sky130_fd_sc_hd__nor2_1 _3896_ (.A(_0683_),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__inv_2 _3897_ (.A(\BitStream_buffer.BS_buffer[80] ),
    .Y(_0686_));
 sky130_fd_sc_hd__o22ai_1 _3898_ (.A1(_0686_),
    .A2(_2697_),
    .B1(_0560_),
    .B2(_2702_),
    .Y(_0687_));
 sky130_fd_sc_hd__a221oi_1 _3899_ (.A1(\BitStream_buffer.BS_buffer[81] ),
    .A2(_2689_),
    .B1(\BitStream_buffer.BS_buffer[82] ),
    .B2(_2693_),
    .C1(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__and4_1 _3900_ (.A(_0678_),
    .B(_0682_),
    .C(_0685_),
    .D(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__or2_1 _3901_ (.A(_0428_),
    .B(_2717_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2_1 _3902_ (.A(_2720_),
    .B(\BitStream_buffer.BS_buffer[93] ),
    .Y(_0691_));
 sky130_fd_sc_hd__nand2_1 _3903_ (.A(_2724_),
    .B(_2714_),
    .Y(_0692_));
 sky130_fd_sc_hd__o2111a_1 _3904_ (.A1(_2737_),
    .A2(_2713_),
    .B1(_0690_),
    .C1(_0691_),
    .D1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__inv_2 _3905_ (.A(_2800_),
    .Y(_0694_));
 sky130_fd_sc_hd__o22ai_1 _3906_ (.A1(_0694_),
    .A2(_2735_),
    .B1(_0568_),
    .B2(_2739_),
    .Y(_0695_));
 sky130_fd_sc_hd__a221oi_1 _3907_ (.A1(\BitStream_buffer.BS_buffer[97] ),
    .A2(_2729_),
    .B1(_2804_),
    .B2(_2732_),
    .C1(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_2746_),
    .B(_2768_),
    .Y(_0697_));
 sky130_fd_sc_hd__nand2_1 _3909_ (.A(_2749_),
    .B(\BitStream_buffer.BS_buffer[83] ),
    .Y(_0698_));
 sky130_fd_sc_hd__or2_1 _3910_ (.A(_0440_),
    .B(_2753_),
    .X(_0699_));
 sky130_fd_sc_hd__o2111a_1 _3911_ (.A1(_0434_),
    .A2(_2744_),
    .B1(_0697_),
    .C1(_0698_),
    .D1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nand2_1 _3912_ (.A(_2761_),
    .B(_2706_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(_2765_),
    .B(_2756_),
    .Y(_0702_));
 sky130_fd_sc_hd__or2_1 _3914_ (.A(_0437_),
    .B(_2771_),
    .X(_0703_));
 sky130_fd_sc_hd__o2111a_1 _3915_ (.A1(_0423_),
    .A2(_2759_),
    .B1(_0701_),
    .C1(_0702_),
    .D1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__and4_1 _3916_ (.A(_0693_),
    .B(_0696_),
    .C(_0700_),
    .D(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__or2_1 _3917_ (.A(_0464_),
    .B(_2784_),
    .X(_0706_));
 sky130_fd_sc_hd__nand2_1 _3918_ (.A(_2787_),
    .B(_2838_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand2_1 _3919_ (.A(_2791_),
    .B(_2781_),
    .Y(_0708_));
 sky130_fd_sc_hd__o2111a_1 _3920_ (.A1(_0445_),
    .A2(_2780_),
    .B1(_0706_),
    .C1(_0707_),
    .D1(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__nand2_1 _3921_ (.A(_2799_),
    .B(\BitStream_buffer.BS_buffer[99] ),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _3922_ (.A(_2803_),
    .B(\BitStream_buffer.BS_buffer[101] ),
    .Y(_0711_));
 sky130_fd_sc_hd__or2_1 _3923_ (.A(_0450_),
    .B(_2808_),
    .X(_0712_));
 sky130_fd_sc_hd__o2111a_1 _3924_ (.A1(_0459_),
    .A2(_2797_),
    .B1(_0710_),
    .C1(_0711_),
    .D1(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__nand2_1 _3925_ (.A(_2815_),
    .B(\BitStream_buffer.BS_buffer[105] ),
    .Y(_0714_));
 sky130_fd_sc_hd__nand2_1 _3926_ (.A(_2819_),
    .B(\BitStream_buffer.BS_buffer[103] ),
    .Y(_0715_));
 sky130_fd_sc_hd__or2_1 _3927_ (.A(_0456_),
    .B(_2824_),
    .X(_0716_));
 sky130_fd_sc_hd__o2111a_1 _3928_ (.A1(_0444_),
    .A2(_2813_),
    .B1(_0714_),
    .C1(_0715_),
    .D1(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__nand2_1 _3929_ (.A(_2831_),
    .B(\BitStream_buffer.BS_buffer[111] ),
    .Y(_0718_));
 sky130_fd_sc_hd__nand2_1 _3930_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[113] ),
    .Y(_0719_));
 sky130_fd_sc_hd__or2_1 _3931_ (.A(_2888_),
    .B(_2841_),
    .X(_0720_));
 sky130_fd_sc_hd__o2111a_1 _3932_ (.A1(_0481_),
    .A2(_2829_),
    .B1(_0718_),
    .C1(_0719_),
    .D1(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__and4_1 _3933_ (.A(_0709_),
    .B(_0713_),
    .C(_0717_),
    .D(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__or2_1 _3934_ (.A(_2883_),
    .B(_2852_),
    .X(_0723_));
 sky130_fd_sc_hd__nand2_1 _3935_ (.A(_2856_),
    .B(\BitStream_buffer.BS_buffer[125] ),
    .Y(_0724_));
 sky130_fd_sc_hd__nand2_1 _3936_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[123] ),
    .Y(_0725_));
 sky130_fd_sc_hd__o2111a_1 _3937_ (.A1(_0476_),
    .A2(_2849_),
    .B1(_0723_),
    .C1(_0724_),
    .D1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__inv_2 _3938_ (.A(\BitStream_buffer.BS_buffer[120] ),
    .Y(_0727_));
 sky130_fd_sc_hd__o22ai_1 _3939_ (.A1(_0727_),
    .A2(_2869_),
    .B1(_0601_),
    .B2(_2872_),
    .Y(_0728_));
 sky130_fd_sc_hd__a221oi_1 _3940_ (.A1(\BitStream_buffer.BS_buffer[121] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[122] ),
    .B2(_2866_),
    .C1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__inv_2 _3941_ (.A(_0400_),
    .Y(_0730_));
 sky130_fd_sc_hd__o22ai_1 _3942_ (.A1(_0730_),
    .A2(_2882_),
    .B1(_0604_),
    .B2(_2885_),
    .Y(_0731_));
 sky130_fd_sc_hd__a221oi_1 _3943_ (.A1(\BitStream_buffer.BS_buffer[1] ),
    .A2(_2876_),
    .B1(_3039_),
    .B2(_2879_),
    .C1(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[117] ),
    .Y(_0733_));
 sky130_fd_sc_hd__or2_1 _3945_ (.A(_0473_),
    .B(_2896_),
    .X(_0734_));
 sky130_fd_sc_hd__or2_1 _3946_ (.A(_2870_),
    .B(_2900_),
    .X(_0735_));
 sky130_fd_sc_hd__o2111a_1 _3947_ (.A1(_2894_),
    .A2(_2890_),
    .B1(_0733_),
    .C1(_0734_),
    .D1(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__and4_1 _3948_ (.A(_0726_),
    .B(_0729_),
    .C(_0732_),
    .D(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__and4_1 _3949_ (.A(_0689_),
    .B(_0705_),
    .C(_0722_),
    .D(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__inv_2 _3950_ (.A(\BitStream_buffer.BS_buffer[40] ),
    .Y(_0739_));
 sky130_fd_sc_hd__o22ai_1 _3951_ (.A1(_0739_),
    .A2(_2909_),
    .B1(_0613_),
    .B2(_2912_),
    .Y(_0740_));
 sky130_fd_sc_hd__o22ai_1 _3952_ (.A1(_0486_),
    .A2(_2916_),
    .B1(_2905_),
    .B2(_2920_),
    .Y(_0741_));
 sky130_fd_sc_hd__a22o_1 _3953_ (.A1(\BitStream_buffer.BS_buffer[41] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[42] ),
    .X(_0742_));
 sky130_fd_sc_hd__a22o_1 _3954_ (.A1(\BitStream_buffer.BS_buffer[35] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[36] ),
    .X(_0743_));
 sky130_fd_sc_hd__or4_1 _3955_ (.A(_0740_),
    .B(_0741_),
    .C(_0742_),
    .D(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__o22ai_1 _3956_ (.A1(_2975_),
    .A2(_2941_),
    .B1(_0619_),
    .B2(_2945_),
    .Y(_0745_));
 sky130_fd_sc_hd__a221oi_1 _3957_ (.A1(\BitStream_buffer.BS_buffer[47] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[48] ),
    .B2(_2938_),
    .C1(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__o22ai_1 _3958_ (.A1(_2942_),
    .A2(_2955_),
    .B1(_0622_),
    .B2(_2959_),
    .Y(_0747_));
 sky130_fd_sc_hd__a221oi_1 _3959_ (.A1(\BitStream_buffer.BS_buffer[43] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[44] ),
    .B2(_2952_),
    .C1(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand3b_1 _3960_ (.A_N(_0744_),
    .B(_0746_),
    .C(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__inv_2 _3961_ (.A(\BitStream_buffer.BS_buffer[56] ),
    .Y(_0750_));
 sky130_fd_sc_hd__o22ai_1 _3962_ (.A1(_0750_),
    .A2(_2967_),
    .B1(_0626_),
    .B2(_2970_),
    .Y(_0751_));
 sky130_fd_sc_hd__o22ai_1 _3963_ (.A1(_0499_),
    .A2(_2974_),
    .B1(_2963_),
    .B2(_2977_),
    .Y(_0752_));
 sky130_fd_sc_hd__a22o_1 _3964_ (.A1(\BitStream_buffer.BS_buffer[57] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[58] ),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_1 _3965_ (.A1(\BitStream_buffer.BS_buffer[51] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[52] ),
    .X(_0754_));
 sky130_fd_sc_hd__or4_1 _3966_ (.A(_0751_),
    .B(_0752_),
    .C(_0753_),
    .D(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__o22ai_1 _3967_ (.A1(_3009_),
    .A2(_2998_),
    .B1(_0632_),
    .B2(_3001_),
    .Y(_0756_));
 sky130_fd_sc_hd__a221oi_1 _3968_ (.A1(\BitStream_buffer.BS_buffer[59] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[60] ),
    .B2(_2995_),
    .C1(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__a2bb2o_1 _3969_ (.A1_N(_2652_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[66] ),
    .B2(_3014_),
    .X(_0758_));
 sky130_fd_sc_hd__a221oi_1 _3970_ (.A1(\BitStream_buffer.BS_buffer[63] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[64] ),
    .B2(_3008_),
    .C1(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__nand3b_1 _3971_ (.A_N(_0755_),
    .B(_0757_),
    .C(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__inv_2 _3972_ (.A(\BitStream_buffer.BS_buffer[4] ),
    .Y(_0761_));
 sky130_fd_sc_hd__nor2_1 _3973_ (.A(_0761_),
    .B(_3022_),
    .Y(_0762_));
 sky130_fd_sc_hd__o22ai_1 _3974_ (.A1(_3063_),
    .A2(_3026_),
    .B1(_0640_),
    .B2(_3030_),
    .Y(_0763_));
 sky130_fd_sc_hd__a22o_1 _3975_ (.A1(\BitStream_buffer.BS_buffer[7] ),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_0330_),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _3976_ (.A1(_3037_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_0516_),
    .X(_0765_));
 sky130_fd_sc_hd__or4_1 _3977_ (.A(_0762_),
    .B(_0763_),
    .C(_0764_),
    .D(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__a22o_1 _3978_ (.A1(\BitStream_buffer.BS_buffer[15] ),
    .A2(_3048_),
    .B1(_3050_),
    .B2(_0363_),
    .X(_0767_));
 sky130_fd_sc_hd__o22ai_1 _3979_ (.A1(_0373_),
    .A2(_3055_),
    .B1(_0646_),
    .B2(_3058_),
    .Y(_0768_));
 sky130_fd_sc_hd__o22ai_1 _3980_ (.A1(_3056_),
    .A2(_3062_),
    .B1(_0648_),
    .B2(_0323_),
    .Y(_0769_));
 sky130_fd_sc_hd__clkbuf_4 _3981_ (.A(\BitStream_buffer.BS_buffer[12] ),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _3982_ (.A1(_0770_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0650_),
    .X(_0771_));
 sky130_fd_sc_hd__or4_1 _3983_ (.A(_0767_),
    .B(_0768_),
    .C(_0769_),
    .D(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__nor2_1 _3984_ (.A(_0766_),
    .B(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__o22ai_1 _3985_ (.A1(_0388_),
    .A2(_0344_),
    .B1(_0654_),
    .B2(_0347_),
    .Y(_0774_));
 sky130_fd_sc_hd__a221oi_1 _3986_ (.A1(\BitStream_buffer.BS_buffer[27] ),
    .A2(_0337_),
    .B1(\BitStream_buffer.BS_buffer[28] ),
    .B2(_0341_),
    .C1(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__o22ai_1 _3987_ (.A1(_0345_),
    .A2(_0357_),
    .B1(_0657_),
    .B2(_0360_),
    .Y(_0776_));
 sky130_fd_sc_hd__a221oi_1 _3988_ (.A1(\BitStream_buffer.BS_buffer[23] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[24] ),
    .B2(_0354_),
    .C1(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__o22ai_1 _3989_ (.A1(_0358_),
    .A2(_0372_),
    .B1(_0660_),
    .B2(_0375_),
    .Y(_0778_));
 sky130_fd_sc_hd__a221oi_1 _3990_ (.A1(\BitStream_buffer.BS_buffer[19] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[20] ),
    .B2(_0369_),
    .C1(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__o22ai_1 _3991_ (.A1(_2917_),
    .A2(_0386_),
    .B1(_0663_),
    .B2(_0390_),
    .Y(_0780_));
 sky130_fd_sc_hd__a221oi_1 _3992_ (.A1(\BitStream_buffer.BS_buffer[32] ),
    .A2(_0382_),
    .B1(\BitStream_buffer.BS_buffer[31] ),
    .B2(_0379_),
    .C1(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__and4_1 _3993_ (.A(_0775_),
    .B(_0777_),
    .C(_0779_),
    .D(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__nand2_1 _3994_ (.A(_0773_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__nor3_1 _3995_ (.A(_0749_),
    .B(_0760_),
    .C(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_0399_),
    .B(_3044_),
    .Y(_0785_));
 sky130_fd_sc_hd__nand3_1 _3997_ (.A(_0738_),
    .B(_0784_),
    .C(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__inv_2 _3998_ (.A(\BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_0787_));
 sky130_fd_sc_hd__a21oi_1 _3999_ (.A1(_0787_),
    .A2(_0672_),
    .B1(_0675_),
    .Y(_0788_));
 sky130_fd_sc_hd__o21a_1 _4000_ (.A1(_2599_),
    .A2(_0786_),
    .B1(_0788_),
    .X(_0318_));
 sky130_fd_sc_hd__o22ai_1 _4001_ (.A1(_2694_),
    .A2(_2630_),
    .B1(_2698_),
    .B2(_2637_),
    .Y(_0789_));
 sky130_fd_sc_hd__a221oi_1 _4002_ (.A1(\BitStream_buffer.BS_buffer[78] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[79] ),
    .B2(_2624_),
    .C1(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nand2_1 _4003_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[70] ),
    .Y(_0791_));
 sky130_fd_sc_hd__or2_1 _4004_ (.A(_2664_),
    .B(_2656_),
    .X(_0792_));
 sky130_fd_sc_hd__or2_1 _4005_ (.A(_0556_),
    .B(_2661_),
    .X(_0793_));
 sky130_fd_sc_hd__o2111a_1 _4006_ (.A1(_2671_),
    .A2(_2646_),
    .B1(_0791_),
    .C1(_0792_),
    .D1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__o22ai_1 _4007_ (.A1(_2625_),
    .A2(_2670_),
    .B1(_2631_),
    .B2(_2675_),
    .Y(_0795_));
 sky130_fd_sc_hd__a22o_1 _4008_ (.A1(\BitStream_buffer.BS_buffer[74] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[75] ),
    .X(_0796_));
 sky130_fd_sc_hd__nor2_1 _4009_ (.A(_0795_),
    .B(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__o22ai_1 _4010_ (.A1(_2742_),
    .A2(_2697_),
    .B1(_0686_),
    .B2(_2702_),
    .Y(_0798_));
 sky130_fd_sc_hd__a221oi_1 _4011_ (.A1(\BitStream_buffer.BS_buffer[82] ),
    .A2(_2689_),
    .B1(\BitStream_buffer.BS_buffer[83] ),
    .B2(_2693_),
    .C1(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__and4_1 _4012_ (.A(_0790_),
    .B(_0794_),
    .C(_0797_),
    .D(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__or2_1 _4013_ (.A(_0568_),
    .B(_2717_),
    .X(_0801_));
 sky130_fd_sc_hd__nand2_1 _4014_ (.A(_2720_),
    .B(\BitStream_buffer.BS_buffer[94] ),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _4015_ (.A(_2724_),
    .B(_2736_),
    .Y(_0803_));
 sky130_fd_sc_hd__o2111a_1 _4016_ (.A1(_2733_),
    .A2(_2713_),
    .B1(_0801_),
    .C1(_0802_),
    .D1(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__o22ai_1 _4017_ (.A1(_2806_),
    .A2(_2735_),
    .B1(_0694_),
    .B2(_2739_),
    .Y(_0805_));
 sky130_fd_sc_hd__a221oi_1 _4018_ (.A1(_2804_),
    .A2(_2729_),
    .B1(\BitStream_buffer.BS_buffer[99] ),
    .B2(_2732_),
    .C1(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(_2746_),
    .B(_2762_),
    .Y(_0807_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_2749_),
    .B(_2766_),
    .Y(_0808_));
 sky130_fd_sc_hd__or2_1 _4021_ (.A(_2757_),
    .B(_2753_),
    .X(_0809_));
 sky130_fd_sc_hd__o2111a_1 _4022_ (.A1(_2769_),
    .A2(_2744_),
    .B1(_0807_),
    .C1(_0808_),
    .D1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_1 _4023_ (.A(_2761_),
    .B(_2721_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _4024_ (.A(_2765_),
    .B(_2725_),
    .Y(_0812_));
 sky130_fd_sc_hd__or2_1 _4025_ (.A(_2707_),
    .B(_2771_),
    .X(_0813_));
 sky130_fd_sc_hd__o2111a_1 _4026_ (.A1(_2715_),
    .A2(_2759_),
    .B1(_0811_),
    .C1(_0812_),
    .D1(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__and4_1 _4027_ (.A(_0804_),
    .B(_0806_),
    .C(_0810_),
    .D(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__or2_1 _4028_ (.A(_2827_),
    .B(_2784_),
    .X(_0816_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(_2787_),
    .B(_2836_),
    .Y(_0817_));
 sky130_fd_sc_hd__nand2_1 _4030_ (.A(_2791_),
    .B(_2832_),
    .Y(_0818_));
 sky130_fd_sc_hd__o2111a_1 _4031_ (.A1(_2839_),
    .A2(_2780_),
    .B1(_0816_),
    .C1(_0817_),
    .D1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__nand2_1 _4032_ (.A(_2799_),
    .B(_2820_),
    .Y(_0820_));
 sky130_fd_sc_hd__nand2_1 _4033_ (.A(_2803_),
    .B(_2816_),
    .Y(_0821_));
 sky130_fd_sc_hd__or2_1 _4034_ (.A(_2822_),
    .B(_2808_),
    .X(_0822_));
 sky130_fd_sc_hd__o2111a_1 _4035_ (.A1(_2811_),
    .A2(_2797_),
    .B1(_0820_),
    .C1(_0821_),
    .D1(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_1 _4036_ (.A(_2815_),
    .B(_2788_),
    .Y(_0824_));
 sky130_fd_sc_hd__nand2_1 _4037_ (.A(_2819_),
    .B(_2792_),
    .Y(_0825_));
 sky130_fd_sc_hd__or2_1 _4038_ (.A(_2775_),
    .B(_2824_),
    .X(_0826_));
 sky130_fd_sc_hd__o2111a_1 _4039_ (.A1(_2782_),
    .A2(_2813_),
    .B1(_0824_),
    .C1(_0825_),
    .D1(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__nand2_1 _4040_ (.A(_2831_),
    .B(\BitStream_buffer.BS_buffer[112] ),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _4041_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[114] ),
    .Y(_0829_));
 sky130_fd_sc_hd__or2_1 _4042_ (.A(_2898_),
    .B(_2841_),
    .X(_0830_));
 sky130_fd_sc_hd__o2111a_1 _4043_ (.A1(_2894_),
    .A2(_2829_),
    .B1(_0828_),
    .C1(_0829_),
    .D1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__and4_1 _4044_ (.A(_0819_),
    .B(_0823_),
    .C(_0827_),
    .D(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__or2_1 _4045_ (.A(_2880_),
    .B(_2852_),
    .X(_0833_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(_2856_),
    .B(\BitStream_buffer.BS_buffer[126] ),
    .Y(_0834_));
 sky130_fd_sc_hd__nand2_1 _4047_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[124] ),
    .Y(_0835_));
 sky130_fd_sc_hd__o2111a_1 _4048_ (.A1(_0604_),
    .A2(_2849_),
    .B1(_0833_),
    .C1(_0834_),
    .D1(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__o22ai_1 _4049_ (.A1(_2850_),
    .A2(_2869_),
    .B1(_0727_),
    .B2(_2872_),
    .Y(_0837_));
 sky130_fd_sc_hd__a221oi_1 _4050_ (.A1(\BitStream_buffer.BS_buffer[122] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[123] ),
    .B2(_2866_),
    .C1(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__o22ai_1 _4051_ (.A1(_3018_),
    .A2(_2882_),
    .B1(_0730_),
    .B2(_2885_),
    .Y(_0839_));
 sky130_fd_sc_hd__a221oi_1 _4052_ (.A1(_3039_),
    .A2(_2876_),
    .B1(_3044_),
    .B2(_2879_),
    .C1(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__nand2_1 _4053_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[118] ),
    .Y(_0841_));
 sky130_fd_sc_hd__or2_1 _4054_ (.A(_0601_),
    .B(_2896_),
    .X(_0842_));
 sky130_fd_sc_hd__or2_1 _4055_ (.A(_2867_),
    .B(_2900_),
    .X(_0843_));
 sky130_fd_sc_hd__o2111a_1 _4056_ (.A1(_2870_),
    .A2(_2890_),
    .B1(_0841_),
    .C1(_0842_),
    .D1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__and4_1 _4057_ (.A(_0836_),
    .B(_0838_),
    .C(_0840_),
    .D(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__and4_1 _4058_ (.A(_0800_),
    .B(_0815_),
    .C(_0832_),
    .D(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__inv_2 _4059_ (.A(\BitStream_buffer.BS_buffer[41] ),
    .Y(_0847_));
 sky130_fd_sc_hd__o22ai_1 _4060_ (.A1(_0847_),
    .A2(_2909_),
    .B1(_0739_),
    .B2(_2912_),
    .Y(_0848_));
 sky130_fd_sc_hd__o22ai_1 _4061_ (.A1(_0613_),
    .A2(_2916_),
    .B1(_0486_),
    .B2(_2920_),
    .Y(_0849_));
 sky130_fd_sc_hd__a22o_1 _4062_ (.A1(\BitStream_buffer.BS_buffer[42] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[43] ),
    .X(_0850_));
 sky130_fd_sc_hd__a22o_1 _4063_ (.A1(\BitStream_buffer.BS_buffer[36] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[37] ),
    .X(_0851_));
 sky130_fd_sc_hd__or4_1 _4064_ (.A(_0848_),
    .B(_0849_),
    .C(_0850_),
    .D(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__o22ai_1 _4065_ (.A1(_2972_),
    .A2(_2941_),
    .B1(_2975_),
    .B2(_2945_),
    .Y(_0853_));
 sky130_fd_sc_hd__a221oi_1 _4066_ (.A1(\BitStream_buffer.BS_buffer[48] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[49] ),
    .B2(_2938_),
    .C1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__o22ai_1 _4067_ (.A1(_2939_),
    .A2(_2955_),
    .B1(_2942_),
    .B2(_2959_),
    .Y(_0855_));
 sky130_fd_sc_hd__a221oi_1 _4068_ (.A1(\BitStream_buffer.BS_buffer[44] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[45] ),
    .B2(_2952_),
    .C1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand3b_1 _4069_ (.A_N(_0852_),
    .B(_0854_),
    .C(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__inv_2 _4070_ (.A(\BitStream_buffer.BS_buffer[57] ),
    .Y(_0858_));
 sky130_fd_sc_hd__o22ai_1 _4071_ (.A1(_0858_),
    .A2(_2967_),
    .B1(_0750_),
    .B2(_2970_),
    .Y(_0859_));
 sky130_fd_sc_hd__o22ai_1 _4072_ (.A1(_0626_),
    .A2(_2974_),
    .B1(_0499_),
    .B2(_2977_),
    .Y(_0860_));
 sky130_fd_sc_hd__a22o_1 _4073_ (.A1(\BitStream_buffer.BS_buffer[58] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[59] ),
    .X(_0861_));
 sky130_fd_sc_hd__a22o_1 _4074_ (.A1(\BitStream_buffer.BS_buffer[52] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[53] ),
    .X(_0862_));
 sky130_fd_sc_hd__or4_1 _4075_ (.A(_0859_),
    .B(_0860_),
    .C(_0861_),
    .D(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__o22ai_1 _4076_ (.A1(_0508_),
    .A2(_2998_),
    .B1(_3009_),
    .B2(_3001_),
    .Y(_0864_));
 sky130_fd_sc_hd__a221oi_1 _4077_ (.A1(\BitStream_buffer.BS_buffer[60] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[61] ),
    .B2(_2995_),
    .C1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__a2bb2o_1 _4078_ (.A1_N(_0411_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[67] ),
    .B2(_3014_),
    .X(_0866_));
 sky130_fd_sc_hd__a221oi_1 _4079_ (.A1(\BitStream_buffer.BS_buffer[64] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[65] ),
    .B2(_3008_),
    .C1(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand3b_1 _4080_ (.A_N(_0863_),
    .B(_0865_),
    .C(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__inv_2 _4081_ (.A(\BitStream_buffer.BS_buffer[5] ),
    .Y(_0869_));
 sky130_fd_sc_hd__nor2_1 _4082_ (.A(_0869_),
    .B(_3022_),
    .Y(_0870_));
 sky130_fd_sc_hd__o22ai_1 _4083_ (.A1(_3060_),
    .A2(_3026_),
    .B1(_3063_),
    .B2(_3030_),
    .Y(_0871_));
 sky130_fd_sc_hd__a22o_1 _4084_ (.A1(_0330_),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_0325_),
    .X(_0872_));
 sky130_fd_sc_hd__a22o_1 _4085_ (.A1(_0516_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(\BitStream_buffer.BS_buffer[7] ),
    .X(_0873_));
 sky130_fd_sc_hd__or4_1 _4086_ (.A(_0870_),
    .B(_0871_),
    .C(_0872_),
    .D(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__a22o_1 _4087_ (.A1(_0363_),
    .A2(_3048_),
    .B1(_3050_),
    .B2(_0366_),
    .X(_0875_));
 sky130_fd_sc_hd__o22ai_1 _4088_ (.A1(_0370_),
    .A2(_3055_),
    .B1(_0373_),
    .B2(_3058_),
    .Y(_0876_));
 sky130_fd_sc_hd__o22ai_1 _4089_ (.A1(_3053_),
    .A2(_3062_),
    .B1(_3056_),
    .B2(_0323_),
    .Y(_0877_));
 sky130_fd_sc_hd__a22o_1 _4090_ (.A1(_3051_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0770_),
    .X(_0878_));
 sky130_fd_sc_hd__or4_1 _4091_ (.A(_0875_),
    .B(_0876_),
    .C(_0877_),
    .D(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_1 _4092_ (.A(_0874_),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__o22ai_1 _4093_ (.A1(_0384_),
    .A2(_0344_),
    .B1(_0388_),
    .B2(_0347_),
    .Y(_0881_));
 sky130_fd_sc_hd__a221oi_1 _4094_ (.A1(\BitStream_buffer.BS_buffer[28] ),
    .A2(_0337_),
    .B1(_0380_),
    .B2(_0341_),
    .C1(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__o22ai_1 _4095_ (.A1(_0342_),
    .A2(_0357_),
    .B1(_0345_),
    .B2(_0360_),
    .Y(_0883_));
 sky130_fd_sc_hd__a221oi_1 _4096_ (.A1(\BitStream_buffer.BS_buffer[24] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[25] ),
    .B2(_0354_),
    .C1(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__o22ai_1 _4097_ (.A1(_0355_),
    .A2(_0372_),
    .B1(_0358_),
    .B2(_0375_),
    .Y(_0885_));
 sky130_fd_sc_hd__a221oi_1 _4098_ (.A1(\BitStream_buffer.BS_buffer[20] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[21] ),
    .B2(_0369_),
    .C1(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__o22ai_1 _4099_ (.A1(_2914_),
    .A2(_0386_),
    .B1(_2917_),
    .B2(_0390_),
    .Y(_0887_));
 sky130_fd_sc_hd__a221oi_2 _4100_ (.A1(\BitStream_buffer.BS_buffer[32] ),
    .A2(_0379_),
    .B1(\BitStream_buffer.BS_buffer[33] ),
    .B2(_0383_),
    .C1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__and4_1 _4101_ (.A(_0882_),
    .B(_0884_),
    .C(_0886_),
    .D(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__nand2_1 _4102_ (.A(_0880_),
    .B(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__nor3_1 _4103_ (.A(_0857_),
    .B(_0868_),
    .C(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_1 _4104_ (.A(_0399_),
    .B(_0518_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand3_1 _4105_ (.A(_0846_),
    .B(_0891_),
    .C(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__inv_4 _4106_ (.A(\BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_0894_));
 sky130_fd_sc_hd__a21oi_1 _4107_ (.A1(_0894_),
    .A2(_0672_),
    .B1(_0675_),
    .Y(_0895_));
 sky130_fd_sc_hd__o21a_1 _4108_ (.A1(_2599_),
    .A2(_0893_),
    .B1(_0895_),
    .X(_0317_));
 sky130_fd_sc_hd__o22ai_1 _4109_ (.A1(_0419_),
    .A2(_2630_),
    .B1(_2694_),
    .B2(_2637_),
    .Y(_0896_));
 sky130_fd_sc_hd__a221oi_1 _4110_ (.A1(\BitStream_buffer.BS_buffer[79] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[80] ),
    .B2(_2624_),
    .C1(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2_1 _4111_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[71] ),
    .Y(_0898_));
 sky130_fd_sc_hd__or2_1 _4112_ (.A(_0415_),
    .B(_2656_),
    .X(_0899_));
 sky130_fd_sc_hd__or2_1 _4113_ (.A(_2631_),
    .B(_2661_),
    .X(_0900_));
 sky130_fd_sc_hd__o2111a_1 _4114_ (.A1(_2664_),
    .A2(_2646_),
    .B1(_0898_),
    .C1(_0899_),
    .D1(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__o22ai_1 _4115_ (.A1(_0407_),
    .A2(_2670_),
    .B1(_2625_),
    .B2(_2675_),
    .Y(_0902_));
 sky130_fd_sc_hd__a22o_1 _4116_ (.A1(\BitStream_buffer.BS_buffer[75] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[76] ),
    .X(_0903_));
 sky130_fd_sc_hd__nor2_1 _4117_ (.A(_0902_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__o22ai_1 _4118_ (.A1(_0431_),
    .A2(_2697_),
    .B1(_2742_),
    .B2(_2702_),
    .Y(_0905_));
 sky130_fd_sc_hd__a221oi_1 _4119_ (.A1(\BitStream_buffer.BS_buffer[83] ),
    .A2(_2689_),
    .B1(_2766_),
    .B2(_2693_),
    .C1(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__and4_1 _4120_ (.A(_0897_),
    .B(_0901_),
    .C(_0904_),
    .D(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__or2_1 _4121_ (.A(_0694_),
    .B(_2717_),
    .X(_0908_));
 sky130_fd_sc_hd__nand2_1 _4122_ (.A(_2720_),
    .B(\BitStream_buffer.BS_buffer[95] ),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_1 _4123_ (.A(_2724_),
    .B(\BitStream_buffer.BS_buffer[93] ),
    .Y(_0910_));
 sky130_fd_sc_hd__o2111a_1 _4124_ (.A1(_0428_),
    .A2(_2713_),
    .B1(_0908_),
    .C1(_0909_),
    .D1(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__o22ai_1 _4125_ (.A1(_0453_),
    .A2(_2735_),
    .B1(_2806_),
    .B2(_2739_),
    .Y(_0912_));
 sky130_fd_sc_hd__a221oi_1 _4126_ (.A1(\BitStream_buffer.BS_buffer[99] ),
    .A2(_2729_),
    .B1(_2820_),
    .B2(_2732_),
    .C1(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__nand2_1 _4127_ (.A(_2746_),
    .B(_2756_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(_2749_),
    .B(_2768_),
    .Y(_0915_));
 sky130_fd_sc_hd__or2_1 _4129_ (.A(_0437_),
    .B(_2753_),
    .X(_0916_));
 sky130_fd_sc_hd__o2111a_1 _4130_ (.A1(_0440_),
    .A2(_2744_),
    .B1(_0914_),
    .C1(_0915_),
    .D1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_1 _4131_ (.A(_2761_),
    .B(_2714_),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _4132_ (.A(_2765_),
    .B(_2706_),
    .Y(_0919_));
 sky130_fd_sc_hd__or2_1 _4133_ (.A(_0423_),
    .B(_2771_),
    .X(_0920_));
 sky130_fd_sc_hd__o2111a_1 _4134_ (.A1(_2737_),
    .A2(_2759_),
    .B1(_0918_),
    .C1(_0919_),
    .D1(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__and4_1 _4135_ (.A(_0911_),
    .B(_0913_),
    .C(_0917_),
    .D(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__or2_1 _4136_ (.A(_2888_),
    .B(_2784_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _4137_ (.A(_2787_),
    .B(\BitStream_buffer.BS_buffer[111] ),
    .Y(_0924_));
 sky130_fd_sc_hd__nand2_1 _4138_ (.A(_2791_),
    .B(_2838_),
    .Y(_0925_));
 sky130_fd_sc_hd__o2111a_1 _4139_ (.A1(_0464_),
    .A2(_2780_),
    .B1(_0923_),
    .C1(_0924_),
    .D1(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__nand2_1 _4140_ (.A(_2799_),
    .B(\BitStream_buffer.BS_buffer[101] ),
    .Y(_0927_));
 sky130_fd_sc_hd__nand2_1 _4141_ (.A(_2803_),
    .B(\BitStream_buffer.BS_buffer[103] ),
    .Y(_0928_));
 sky130_fd_sc_hd__or2_1 _4142_ (.A(_0459_),
    .B(_2808_),
    .X(_0929_));
 sky130_fd_sc_hd__o2111a_1 _4143_ (.A1(_0456_),
    .A2(_2797_),
    .B1(_0927_),
    .C1(_0928_),
    .D1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__nand2_1 _4144_ (.A(_2815_),
    .B(_2781_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _4145_ (.A(_2819_),
    .B(\BitStream_buffer.BS_buffer[105] ),
    .Y(_0932_));
 sky130_fd_sc_hd__or2_1 _4146_ (.A(_0444_),
    .B(_2824_),
    .X(_0933_));
 sky130_fd_sc_hd__o2111a_1 _4147_ (.A1(_0445_),
    .A2(_2813_),
    .B1(_0931_),
    .C1(_0932_),
    .D1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__nand2_1 _4148_ (.A(_2831_),
    .B(\BitStream_buffer.BS_buffer[113] ),
    .Y(_0935_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[115] ),
    .Y(_0936_));
 sky130_fd_sc_hd__or2_1 _4150_ (.A(_0481_),
    .B(_2841_),
    .X(_0937_));
 sky130_fd_sc_hd__o2111a_1 _4151_ (.A1(_2870_),
    .A2(_2829_),
    .B1(_0935_),
    .C1(_0936_),
    .D1(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__and4_1 _4152_ (.A(_0926_),
    .B(_0930_),
    .C(_0934_),
    .D(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__or2_1 _4153_ (.A(_0476_),
    .B(_2852_),
    .X(_0940_));
 sky130_fd_sc_hd__nand2_1 _4154_ (.A(_2856_),
    .B(\BitStream_buffer.BS_buffer[127] ),
    .Y(_0941_));
 sky130_fd_sc_hd__nand2_1 _4155_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[125] ),
    .Y(_0942_));
 sky130_fd_sc_hd__o2111a_1 _4156_ (.A1(_0730_),
    .A2(_2849_),
    .B1(_0940_),
    .C1(_0941_),
    .D1(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__o22ai_1 _4157_ (.A1(_0468_),
    .A2(_2869_),
    .B1(_2850_),
    .B2(_2872_),
    .Y(_0944_));
 sky130_fd_sc_hd__a221oi_1 _4158_ (.A1(\BitStream_buffer.BS_buffer[123] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[124] ),
    .B2(_2866_),
    .C1(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__o22ai_1 _4159_ (.A1(_0512_),
    .A2(_2882_),
    .B1(_3018_),
    .B2(_2885_),
    .Y(_0946_));
 sky130_fd_sc_hd__a221oi_1 _4160_ (.A1(_3044_),
    .A2(_2876_),
    .B1(_0518_),
    .B2(_2879_),
    .C1(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _4161_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[119] ),
    .Y(_0948_));
 sky130_fd_sc_hd__or2_1 _4162_ (.A(_0727_),
    .B(_2896_),
    .X(_0949_));
 sky130_fd_sc_hd__or2_1 _4163_ (.A(_0473_),
    .B(_2900_),
    .X(_0950_));
 sky130_fd_sc_hd__o2111a_1 _4164_ (.A1(_2867_),
    .A2(_2890_),
    .B1(_0948_),
    .C1(_0949_),
    .D1(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__and4_1 _4165_ (.A(_0943_),
    .B(_0945_),
    .C(_0947_),
    .D(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__and4_1 _4166_ (.A(_0907_),
    .B(_0922_),
    .C(_0939_),
    .D(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__o22ai_1 _4167_ (.A1(_2956_),
    .A2(_2909_),
    .B1(_0847_),
    .B2(_2912_),
    .Y(_0954_));
 sky130_fd_sc_hd__o22ai_1 _4168_ (.A1(_0739_),
    .A2(_2916_),
    .B1(_0613_),
    .B2(_2920_),
    .Y(_0955_));
 sky130_fd_sc_hd__a22o_1 _4169_ (.A1(\BitStream_buffer.BS_buffer[43] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[44] ),
    .X(_0956_));
 sky130_fd_sc_hd__a22o_1 _4170_ (.A1(\BitStream_buffer.BS_buffer[37] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[38] ),
    .X(_0957_));
 sky130_fd_sc_hd__or4_1 _4171_ (.A(_0954_),
    .B(_0955_),
    .C(_0956_),
    .D(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__o22ai_1 _4172_ (.A1(_2968_),
    .A2(_2941_),
    .B1(_2972_),
    .B2(_2945_),
    .Y(_0959_));
 sky130_fd_sc_hd__a221oi_2 _4173_ (.A1(\BitStream_buffer.BS_buffer[49] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[50] ),
    .B2(_2938_),
    .C1(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__o22ai_1 _4174_ (.A1(_0492_),
    .A2(_2955_),
    .B1(_2939_),
    .B2(_2959_),
    .Y(_0961_));
 sky130_fd_sc_hd__a221oi_1 _4175_ (.A1(\BitStream_buffer.BS_buffer[45] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[46] ),
    .B2(_2952_),
    .C1(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__nand3b_1 _4176_ (.A_N(_0958_),
    .B(_0960_),
    .C(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__o22ai_1 _4177_ (.A1(_2999_),
    .A2(_2967_),
    .B1(_0858_),
    .B2(_2970_),
    .Y(_0964_));
 sky130_fd_sc_hd__o22ai_1 _4178_ (.A1(_0750_),
    .A2(_2974_),
    .B1(_0626_),
    .B2(_2977_),
    .Y(_0965_));
 sky130_fd_sc_hd__a22o_1 _4179_ (.A1(\BitStream_buffer.BS_buffer[59] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[60] ),
    .X(_0966_));
 sky130_fd_sc_hd__a22o_1 _4180_ (.A1(\BitStream_buffer.BS_buffer[53] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[54] ),
    .X(_0967_));
 sky130_fd_sc_hd__or4_1 _4181_ (.A(_0964_),
    .B(_0965_),
    .C(_0966_),
    .D(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__o22ai_1 _4182_ (.A1(_2640_),
    .A2(_2998_),
    .B1(_0508_),
    .B2(_3001_),
    .Y(_0969_));
 sky130_fd_sc_hd__a221oi_1 _4183_ (.A1(\BitStream_buffer.BS_buffer[61] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[62] ),
    .B2(_2995_),
    .C1(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__a2bb2o_1 _4184_ (.A1_N(_2658_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[68] ),
    .B2(_3014_),
    .X(_0971_));
 sky130_fd_sc_hd__a221oi_1 _4185_ (.A1(\BitStream_buffer.BS_buffer[65] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[66] ),
    .B2(_3008_),
    .C1(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__nand3b_1 _4186_ (.A_N(_0968_),
    .B(_0970_),
    .C(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__nor2_1 _4187_ (.A(_3027_),
    .B(_3022_),
    .Y(_0974_));
 sky130_fd_sc_hd__o22ai_1 _4188_ (.A1(_0525_),
    .A2(_3026_),
    .B1(_3060_),
    .B2(_3030_),
    .Y(_0975_));
 sky130_fd_sc_hd__a22o_1 _4189_ (.A1(_0325_),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_0527_),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _4190_ (.A1(\BitStream_buffer.BS_buffer[7] ),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_0330_),
    .X(_0977_));
 sky130_fd_sc_hd__or4_1 _4191_ (.A(_0974_),
    .B(_0975_),
    .C(_0976_),
    .D(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__a22o_1 _4192_ (.A1(_0366_),
    .A2(_3048_),
    .B1(_3050_),
    .B2(\BitStream_buffer.BS_buffer[18] ),
    .X(_0979_));
 sky130_fd_sc_hd__o22ai_1 _4193_ (.A1(_0537_),
    .A2(_3055_),
    .B1(_0370_),
    .B2(_3058_),
    .Y(_0980_));
 sky130_fd_sc_hd__o22ai_1 _4194_ (.A1(_0523_),
    .A2(_3062_),
    .B1(_3053_),
    .B2(_0323_),
    .Y(_0981_));
 sky130_fd_sc_hd__a22o_1 _4195_ (.A1(_0521_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_3051_),
    .X(_0982_));
 sky130_fd_sc_hd__or4_1 _4196_ (.A(_0979_),
    .B(_0980_),
    .C(_0981_),
    .D(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__nor2_1 _4197_ (.A(_0978_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__o22ai_1 _4198_ (.A1(_0540_),
    .A2(_0344_),
    .B1(_0384_),
    .B2(_0347_),
    .Y(_0985_));
 sky130_fd_sc_hd__a221oi_1 _4199_ (.A1(_0380_),
    .A2(_0337_),
    .B1(_0387_),
    .B2(_0341_),
    .C1(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__o22ai_1 _4200_ (.A1(_0531_),
    .A2(_0357_),
    .B1(_0342_),
    .B2(_0360_),
    .Y(_0987_));
 sky130_fd_sc_hd__a221oi_1 _4201_ (.A1(\BitStream_buffer.BS_buffer[25] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[26] ),
    .B2(_0354_),
    .C1(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__o22ai_1 _4202_ (.A1(_0534_),
    .A2(_0372_),
    .B1(_0355_),
    .B2(_0375_),
    .Y(_0989_));
 sky130_fd_sc_hd__a221oi_1 _4203_ (.A1(\BitStream_buffer.BS_buffer[21] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[22] ),
    .B2(_0369_),
    .C1(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__o22ai_1 _4204_ (.A1(_2910_),
    .A2(_0386_),
    .B1(_2914_),
    .B2(_0390_),
    .Y(_0991_));
 sky130_fd_sc_hd__a221oi_1 _4205_ (.A1(\BitStream_buffer.BS_buffer[33] ),
    .A2(_0379_),
    .B1(\BitStream_buffer.BS_buffer[34] ),
    .B2(_0383_),
    .C1(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__and4_1 _4206_ (.A(_0986_),
    .B(_0988_),
    .C(_0990_),
    .D(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__nand2_1 _4207_ (.A(_0984_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__nor3_1 _4208_ (.A(_0963_),
    .B(_0973_),
    .C(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _4209_ (.A(_0399_),
    .B(_3037_),
    .Y(_0996_));
 sky130_fd_sc_hd__nand3_1 _4210_ (.A(_0953_),
    .B(_0995_),
    .C(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__inv_2 _4211_ (.A(\BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_0998_));
 sky130_fd_sc_hd__a21oi_1 _4212_ (.A1(_0998_),
    .A2(_0672_),
    .B1(_0675_),
    .Y(_0999_));
 sky130_fd_sc_hd__o21a_1 _4213_ (.A1(_2599_),
    .A2(_0997_),
    .B1(_0999_),
    .X(_0316_));
 sky130_fd_sc_hd__o22ai_1 _4214_ (.A1(_0560_),
    .A2(_2630_),
    .B1(_0419_),
    .B2(_2637_),
    .Y(_1000_));
 sky130_fd_sc_hd__a221oi_1 _4215_ (.A1(\BitStream_buffer.BS_buffer[80] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[81] ),
    .B2(_2624_),
    .C1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__nand2_1 _4216_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[72] ),
    .Y(_1002_));
 sky130_fd_sc_hd__or2_1 _4217_ (.A(_0556_),
    .B(_2656_),
    .X(_1003_));
 sky130_fd_sc_hd__or2_1 _4218_ (.A(_2625_),
    .B(_2661_),
    .X(_1004_));
 sky130_fd_sc_hd__o2111a_1 _4219_ (.A1(_0415_),
    .A2(_2646_),
    .B1(_1002_),
    .C1(_1003_),
    .D1(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__o22ai_1 _4220_ (.A1(_0549_),
    .A2(_2670_),
    .B1(_0407_),
    .B2(_2675_),
    .Y(_1006_));
 sky130_fd_sc_hd__a22o_1 _4221_ (.A1(\BitStream_buffer.BS_buffer[76] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[77] ),
    .X(_1007_));
 sky130_fd_sc_hd__nor2_1 _4222_ (.A(_1006_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__o22ai_1 _4223_ (.A1(_2751_),
    .A2(_2697_),
    .B1(_0431_),
    .B2(_2702_),
    .Y(_1009_));
 sky130_fd_sc_hd__a221oi_1 _4224_ (.A1(_2766_),
    .A2(_2689_),
    .B1(_2768_),
    .B2(_2693_),
    .C1(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__and4_1 _4225_ (.A(_1001_),
    .B(_1005_),
    .C(_1008_),
    .D(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__or2_1 _4226_ (.A(_2806_),
    .B(_2717_),
    .X(_1012_));
 sky130_fd_sc_hd__nand2_1 _4227_ (.A(_2720_),
    .B(_2800_),
    .Y(_1013_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(_2724_),
    .B(\BitStream_buffer.BS_buffer[94] ),
    .Y(_1014_));
 sky130_fd_sc_hd__o2111a_1 _4229_ (.A1(_0568_),
    .A2(_2713_),
    .B1(_1012_),
    .C1(_1013_),
    .D1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__o22ai_1 _4230_ (.A1(_2795_),
    .A2(_2735_),
    .B1(_0453_),
    .B2(_2739_),
    .Y(_1016_));
 sky130_fd_sc_hd__a221oi_1 _4231_ (.A1(_2820_),
    .A2(_2729_),
    .B1(\BitStream_buffer.BS_buffer[101] ),
    .B2(_2732_),
    .C1(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__nand2_1 _4232_ (.A(_2746_),
    .B(_2725_),
    .Y(_1018_));
 sky130_fd_sc_hd__nand2_1 _4233_ (.A(_2749_),
    .B(_2762_),
    .Y(_1019_));
 sky130_fd_sc_hd__or2_1 _4234_ (.A(_2707_),
    .B(_2753_),
    .X(_1020_));
 sky130_fd_sc_hd__o2111a_1 _4235_ (.A1(_2757_),
    .A2(_2744_),
    .B1(_1018_),
    .C1(_1019_),
    .D1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__nand2_1 _4236_ (.A(_2761_),
    .B(_2736_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2_1 _4237_ (.A(_2765_),
    .B(_2721_),
    .Y(_1023_));
 sky130_fd_sc_hd__or2_1 _4238_ (.A(_2715_),
    .B(_2771_),
    .X(_1024_));
 sky130_fd_sc_hd__o2111a_1 _4239_ (.A1(_2733_),
    .A2(_2759_),
    .B1(_1022_),
    .C1(_1023_),
    .D1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__and4_1 _4240_ (.A(_1015_),
    .B(_1017_),
    .C(_1021_),
    .D(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__or2_1 _4241_ (.A(_2898_),
    .B(_2784_),
    .X(_1027_));
 sky130_fd_sc_hd__nand2_1 _4242_ (.A(_2787_),
    .B(\BitStream_buffer.BS_buffer[112] ),
    .Y(_1028_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(_2791_),
    .B(_2836_),
    .Y(_1029_));
 sky130_fd_sc_hd__o2111a_1 _4244_ (.A1(_2827_),
    .A2(_2780_),
    .B1(_1027_),
    .C1(_1028_),
    .D1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__nand2_1 _4245_ (.A(_2799_),
    .B(_2816_),
    .Y(_1031_));
 sky130_fd_sc_hd__nand2_1 _4246_ (.A(_2803_),
    .B(_2792_),
    .Y(_1032_));
 sky130_fd_sc_hd__or2_1 _4247_ (.A(_2811_),
    .B(_2808_),
    .X(_1033_));
 sky130_fd_sc_hd__o2111a_1 _4248_ (.A1(_2775_),
    .A2(_2797_),
    .B1(_1031_),
    .C1(_1032_),
    .D1(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__nand2_1 _4249_ (.A(_2815_),
    .B(_2832_),
    .Y(_1035_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(_2819_),
    .B(_2788_),
    .Y(_1036_));
 sky130_fd_sc_hd__or2_1 _4251_ (.A(_2782_),
    .B(_2824_),
    .X(_1037_));
 sky130_fd_sc_hd__o2111a_1 _4252_ (.A1(_2839_),
    .A2(_2813_),
    .B1(_1035_),
    .C1(_1036_),
    .D1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(_2831_),
    .B(\BitStream_buffer.BS_buffer[114] ),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _4254_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[116] ),
    .Y(_1040_));
 sky130_fd_sc_hd__or2_1 _4255_ (.A(_2894_),
    .B(_2841_),
    .X(_1041_));
 sky130_fd_sc_hd__o2111a_1 _4256_ (.A1(_2867_),
    .A2(_2829_),
    .B1(_1039_),
    .C1(_1040_),
    .D1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__and4_1 _4257_ (.A(_1030_),
    .B(_1034_),
    .C(_1038_),
    .D(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__or2_1 _4258_ (.A(_0604_),
    .B(_2852_),
    .X(_1044_));
 sky130_fd_sc_hd__nand2_1 _4259_ (.A(_2856_),
    .B(_0400_),
    .Y(_1045_));
 sky130_fd_sc_hd__nand2_1 _4260_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[126] ),
    .Y(_1046_));
 sky130_fd_sc_hd__o2111a_1 _4261_ (.A1(_3018_),
    .A2(_2849_),
    .B1(_1044_),
    .C1(_1045_),
    .D1(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__o22ai_1 _4262_ (.A1(_2845_),
    .A2(_2869_),
    .B1(_0468_),
    .B2(_2872_),
    .Y(_1048_));
 sky130_fd_sc_hd__a221oi_1 _4263_ (.A1(\BitStream_buffer.BS_buffer[124] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[125] ),
    .B2(_2866_),
    .C1(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__o22ai_1 _4264_ (.A1(_0638_),
    .A2(_2882_),
    .B1(_0512_),
    .B2(_2885_),
    .Y(_1050_));
 sky130_fd_sc_hd__a221oi_1 _4265_ (.A1(_0518_),
    .A2(_2876_),
    .B1(_3037_),
    .B2(_2879_),
    .C1(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__nand2_1 _4266_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[120] ),
    .Y(_1052_));
 sky130_fd_sc_hd__or2_1 _4267_ (.A(_2850_),
    .B(_2896_),
    .X(_1053_));
 sky130_fd_sc_hd__or2_1 _4268_ (.A(_0601_),
    .B(_2900_),
    .X(_1054_));
 sky130_fd_sc_hd__o2111a_1 _4269_ (.A1(_0473_),
    .A2(_2890_),
    .B1(_1052_),
    .C1(_1053_),
    .D1(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__and4_1 _4270_ (.A(_1047_),
    .B(_1049_),
    .C(_1051_),
    .D(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__and4_1 _4271_ (.A(_1011_),
    .B(_1026_),
    .C(_1043_),
    .D(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__o22ai_1 _4272_ (.A1(_2953_),
    .A2(_2909_),
    .B1(_2956_),
    .B2(_2912_),
    .Y(_1058_));
 sky130_fd_sc_hd__o22ai_1 _4273_ (.A1(_0847_),
    .A2(_2916_),
    .B1(_0739_),
    .B2(_2920_),
    .Y(_1059_));
 sky130_fd_sc_hd__a22o_1 _4274_ (.A1(\BitStream_buffer.BS_buffer[44] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[45] ),
    .X(_1060_));
 sky130_fd_sc_hd__a22o_1 _4275_ (.A1(\BitStream_buffer.BS_buffer[38] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[39] ),
    .X(_1061_));
 sky130_fd_sc_hd__or4_1 _4276_ (.A(_1058_),
    .B(_1059_),
    .C(_1060_),
    .D(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__o22ai_1 _4277_ (.A1(_2963_),
    .A2(_2941_),
    .B1(_2968_),
    .B2(_2945_),
    .Y(_1063_));
 sky130_fd_sc_hd__a221oi_1 _4278_ (.A1(\BitStream_buffer.BS_buffer[50] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[51] ),
    .B2(_2938_),
    .C1(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__o22ai_1 _4279_ (.A1(_0619_),
    .A2(_2955_),
    .B1(_0492_),
    .B2(_2959_),
    .Y(_1065_));
 sky130_fd_sc_hd__a221oi_1 _4280_ (.A1(\BitStream_buffer.BS_buffer[46] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[47] ),
    .B2(_2952_),
    .C1(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__nand3b_1 _4281_ (.A_N(_1062_),
    .B(_1064_),
    .C(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__o22ai_1 _4282_ (.A1(_2996_),
    .A2(_2967_),
    .B1(_2999_),
    .B2(_2970_),
    .Y(_1068_));
 sky130_fd_sc_hd__o22ai_1 _4283_ (.A1(_0858_),
    .A2(_2974_),
    .B1(_0750_),
    .B2(_2977_),
    .Y(_1069_));
 sky130_fd_sc_hd__a22o_1 _4284_ (.A1(\BitStream_buffer.BS_buffer[60] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[61] ),
    .X(_1070_));
 sky130_fd_sc_hd__a22o_1 _4285_ (.A1(\BitStream_buffer.BS_buffer[54] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[55] ),
    .X(_1071_));
 sky130_fd_sc_hd__or4_1 _4286_ (.A(_1068_),
    .B(_1069_),
    .C(_1070_),
    .D(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__o22ai_1 _4287_ (.A1(_2652_),
    .A2(_2998_),
    .B1(_2640_),
    .B2(_3001_),
    .Y(_1073_));
 sky130_fd_sc_hd__a221oi_1 _4288_ (.A1(\BitStream_buffer.BS_buffer[62] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[63] ),
    .B2(_2995_),
    .C1(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__a2bb2o_1 _4289_ (.A1_N(_2671_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[69] ),
    .B2(_3014_),
    .X(_1075_));
 sky130_fd_sc_hd__a221oi_1 _4290_ (.A1(\BitStream_buffer.BS_buffer[66] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[67] ),
    .B2(_3008_),
    .C1(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__nand3b_1 _4291_ (.A_N(_1072_),
    .B(_1074_),
    .C(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__nor2_1 _4292_ (.A(_3024_),
    .B(_3022_),
    .Y(_1078_));
 sky130_fd_sc_hd__o22ai_1 _4293_ (.A1(_0648_),
    .A2(_3026_),
    .B1(_0525_),
    .B2(_3030_),
    .Y(_1079_));
 sky130_fd_sc_hd__a22o_1 _4294_ (.A1(_0527_),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_0650_),
    .X(_1080_));
 sky130_fd_sc_hd__a22o_1 _4295_ (.A1(_0330_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_0325_),
    .X(_1081_));
 sky130_fd_sc_hd__or4_1 _4296_ (.A(_1078_),
    .B(_1079_),
    .C(_1080_),
    .D(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__a22o_1 _4297_ (.A1(\BitStream_buffer.BS_buffer[18] ),
    .A2(_3048_),
    .B1(_3050_),
    .B2(\BitStream_buffer.BS_buffer[19] ),
    .X(_1083_));
 sky130_fd_sc_hd__o22ai_1 _4298_ (.A1(_0660_),
    .A2(_3055_),
    .B1(_0537_),
    .B2(_3058_),
    .Y(_1084_));
 sky130_fd_sc_hd__o22ai_1 _4299_ (.A1(_0646_),
    .A2(_3062_),
    .B1(_0523_),
    .B2(_0323_),
    .Y(_1085_));
 sky130_fd_sc_hd__a22o_1 _4300_ (.A1(\BitStream_buffer.BS_buffer[15] ),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0521_),
    .X(_1086_));
 sky130_fd_sc_hd__or4_1 _4301_ (.A(_1083_),
    .B(_1084_),
    .C(_1085_),
    .D(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_1 _4302_ (.A(_1082_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__o22ai_1 _4303_ (.A1(_0663_),
    .A2(_0344_),
    .B1(_0540_),
    .B2(_0347_),
    .Y(_1089_));
 sky130_fd_sc_hd__a221oi_1 _4304_ (.A1(_0387_),
    .A2(_0337_),
    .B1(\BitStream_buffer.BS_buffer[31] ),
    .B2(_0341_),
    .C1(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__o22ai_1 _4305_ (.A1(_0654_),
    .A2(_0357_),
    .B1(_0531_),
    .B2(_0360_),
    .Y(_1091_));
 sky130_fd_sc_hd__a221oi_1 _4306_ (.A1(\BitStream_buffer.BS_buffer[26] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[27] ),
    .B2(_0354_),
    .C1(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__o22ai_1 _4307_ (.A1(_0657_),
    .A2(_0372_),
    .B1(_0534_),
    .B2(_0375_),
    .Y(_1093_));
 sky130_fd_sc_hd__a221oi_1 _4308_ (.A1(\BitStream_buffer.BS_buffer[22] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[23] ),
    .B2(_0369_),
    .C1(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__o22ai_1 _4309_ (.A1(_2905_),
    .A2(_0386_),
    .B1(_2910_),
    .B2(_0390_),
    .Y(_1095_));
 sky130_fd_sc_hd__a221oi_1 _4310_ (.A1(\BitStream_buffer.BS_buffer[34] ),
    .A2(_0379_),
    .B1(\BitStream_buffer.BS_buffer[35] ),
    .B2(_0383_),
    .C1(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__and4_1 _4311_ (.A(_1090_),
    .B(_1092_),
    .C(_1094_),
    .D(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_1088_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__nor3_1 _4313_ (.A(_1067_),
    .B(_1077_),
    .C(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_0399_),
    .B(_0516_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand3_1 _4315_ (.A(_1057_),
    .B(_1099_),
    .C(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__inv_2 _4316_ (.A(\BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_1102_));
 sky130_fd_sc_hd__a21oi_1 _4317_ (.A1(_1102_),
    .A2(_0672_),
    .B1(_0674_),
    .Y(_1103_));
 sky130_fd_sc_hd__o21a_1 _4318_ (.A1(_2599_),
    .A2(_1101_),
    .B1(_1103_),
    .X(_0315_));
 sky130_fd_sc_hd__o22ai_1 _4319_ (.A1(_0686_),
    .A2(_2630_),
    .B1(_0560_),
    .B2(_2637_),
    .Y(_1104_));
 sky130_fd_sc_hd__a221oi_1 _4320_ (.A1(\BitStream_buffer.BS_buffer[81] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[82] ),
    .B2(_2624_),
    .C1(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__nand2_1 _4321_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[73] ),
    .Y(_1106_));
 sky130_fd_sc_hd__or2_1 _4322_ (.A(_2631_),
    .B(_2656_),
    .X(_1107_));
 sky130_fd_sc_hd__or2_1 _4323_ (.A(_0407_),
    .B(_2661_),
    .X(_1108_));
 sky130_fd_sc_hd__o2111a_1 _4324_ (.A1(_0556_),
    .A2(_2646_),
    .B1(_1106_),
    .C1(_1107_),
    .D1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__o22ai_1 _4325_ (.A1(_2698_),
    .A2(_2670_),
    .B1(_0549_),
    .B2(_2675_),
    .Y(_1110_));
 sky130_fd_sc_hd__a22o_1 _4326_ (.A1(\BitStream_buffer.BS_buffer[77] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[78] ),
    .X(_1111_));
 sky130_fd_sc_hd__nor2_1 _4327_ (.A(_1110_),
    .B(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__o22ai_1 _4328_ (.A1(_0434_),
    .A2(_2697_),
    .B1(_2751_),
    .B2(_2702_),
    .Y(_1113_));
 sky130_fd_sc_hd__a221oi_1 _4329_ (.A1(_2768_),
    .A2(_2689_),
    .B1(_2762_),
    .B2(_2693_),
    .C1(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__and4_1 _4330_ (.A(_1105_),
    .B(_1109_),
    .C(_1112_),
    .D(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__or2_1 _4331_ (.A(_0453_),
    .B(_2717_),
    .X(_1116_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_2720_),
    .B(\BitStream_buffer.BS_buffer[97] ),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(_2724_),
    .B(\BitStream_buffer.BS_buffer[95] ),
    .Y(_1118_));
 sky130_fd_sc_hd__o2111a_1 _4334_ (.A1(_0694_),
    .A2(_2713_),
    .B1(_1116_),
    .C1(_1117_),
    .D1(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__o22ai_1 _4335_ (.A1(_0450_),
    .A2(_2735_),
    .B1(_2795_),
    .B2(_2739_),
    .Y(_1120_));
 sky130_fd_sc_hd__a221oi_1 _4336_ (.A1(\BitStream_buffer.BS_buffer[101] ),
    .A2(_2729_),
    .B1(_2816_),
    .B2(_2732_),
    .C1(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_2746_),
    .B(_2706_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand2_1 _4338_ (.A(_2749_),
    .B(_2756_),
    .Y(_1123_));
 sky130_fd_sc_hd__or2_1 _4339_ (.A(_0423_),
    .B(_2753_),
    .X(_1124_));
 sky130_fd_sc_hd__o2111a_1 _4340_ (.A1(_0437_),
    .A2(_2744_),
    .B1(_1122_),
    .C1(_1123_),
    .D1(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nand2_1 _4341_ (.A(_2761_),
    .B(\BitStream_buffer.BS_buffer[93] ),
    .Y(_1126_));
 sky130_fd_sc_hd__nand2_1 _4342_ (.A(_2765_),
    .B(_2714_),
    .Y(_1127_));
 sky130_fd_sc_hd__or2_1 _4343_ (.A(_2737_),
    .B(_2771_),
    .X(_1128_));
 sky130_fd_sc_hd__o2111a_1 _4344_ (.A1(_0428_),
    .A2(_2759_),
    .B1(_1126_),
    .C1(_1127_),
    .D1(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__and4_1 _4345_ (.A(_1119_),
    .B(_1121_),
    .C(_1125_),
    .D(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__or2_1 _4346_ (.A(_0481_),
    .B(_2784_),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _4347_ (.A(_2787_),
    .B(\BitStream_buffer.BS_buffer[113] ),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_1 _4348_ (.A(_2791_),
    .B(\BitStream_buffer.BS_buffer[111] ),
    .Y(_1133_));
 sky130_fd_sc_hd__o2111a_1 _4349_ (.A1(_2888_),
    .A2(_2780_),
    .B1(_1131_),
    .C1(_1132_),
    .D1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _4350_ (.A(_2799_),
    .B(\BitStream_buffer.BS_buffer[103] ),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _4351_ (.A(_2803_),
    .B(\BitStream_buffer.BS_buffer[105] ),
    .Y(_1136_));
 sky130_fd_sc_hd__or2_1 _4352_ (.A(_0456_),
    .B(_2808_),
    .X(_1137_));
 sky130_fd_sc_hd__o2111a_1 _4353_ (.A1(_0444_),
    .A2(_2797_),
    .B1(_1135_),
    .C1(_1136_),
    .D1(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_2815_),
    .B(_2838_),
    .Y(_1139_));
 sky130_fd_sc_hd__nand2_1 _4355_ (.A(_2819_),
    .B(_2781_),
    .Y(_1140_));
 sky130_fd_sc_hd__or2_1 _4356_ (.A(_0445_),
    .B(_2824_),
    .X(_1141_));
 sky130_fd_sc_hd__o2111a_1 _4357_ (.A1(_0464_),
    .A2(_2813_),
    .B1(_1139_),
    .C1(_1140_),
    .D1(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__nand2_1 _4358_ (.A(_2831_),
    .B(\BitStream_buffer.BS_buffer[115] ),
    .Y(_1143_));
 sky130_fd_sc_hd__nand2_1 _4359_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[117] ),
    .Y(_1144_));
 sky130_fd_sc_hd__or2_1 _4360_ (.A(_2870_),
    .B(_2841_),
    .X(_1145_));
 sky130_fd_sc_hd__o2111a_1 _4361_ (.A1(_0473_),
    .A2(_2829_),
    .B1(_1143_),
    .C1(_1144_),
    .D1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__and4_1 _4362_ (.A(_1134_),
    .B(_1138_),
    .C(_1142_),
    .D(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__or2_1 _4363_ (.A(_0730_),
    .B(_2852_),
    .X(_1148_));
 sky130_fd_sc_hd__nand2_1 _4364_ (.A(_2856_),
    .B(\BitStream_buffer.BS_buffer[1] ),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[127] ),
    .Y(_1150_));
 sky130_fd_sc_hd__o2111a_1 _4366_ (.A1(_0512_),
    .A2(_2849_),
    .B1(_1148_),
    .C1(_1149_),
    .D1(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__o22ai_1 _4367_ (.A1(_2883_),
    .A2(_2869_),
    .B1(_2845_),
    .B2(_2872_),
    .Y(_1152_));
 sky130_fd_sc_hd__a221oi_1 _4368_ (.A1(\BitStream_buffer.BS_buffer[125] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[126] ),
    .B2(_2866_),
    .C1(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__o22ai_1 _4369_ (.A1(_0761_),
    .A2(_2882_),
    .B1(_0638_),
    .B2(_2885_),
    .Y(_1154_));
 sky130_fd_sc_hd__a221oi_1 _4370_ (.A1(_3037_),
    .A2(_2876_),
    .B1(_0516_),
    .B2(_2879_),
    .C1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__nand2_1 _4371_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[121] ),
    .Y(_1156_));
 sky130_fd_sc_hd__or2_1 _4372_ (.A(_0468_),
    .B(_2896_),
    .X(_1157_));
 sky130_fd_sc_hd__or2_1 _4373_ (.A(_0727_),
    .B(_2900_),
    .X(_1158_));
 sky130_fd_sc_hd__o2111a_1 _4374_ (.A1(_0601_),
    .A2(_2890_),
    .B1(_1156_),
    .C1(_1157_),
    .D1(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__and4_1 _4375_ (.A(_1151_),
    .B(_1153_),
    .C(_1155_),
    .D(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__and4_1 _4376_ (.A(_1115_),
    .B(_1130_),
    .C(_1147_),
    .D(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__o22ai_1 _4377_ (.A1(_0495_),
    .A2(_2909_),
    .B1(_2953_),
    .B2(_2912_),
    .Y(_1162_));
 sky130_fd_sc_hd__o22ai_1 _4378_ (.A1(_2956_),
    .A2(_2916_),
    .B1(_0847_),
    .B2(_2920_),
    .Y(_1163_));
 sky130_fd_sc_hd__a22o_1 _4379_ (.A1(\BitStream_buffer.BS_buffer[45] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[46] ),
    .X(_1164_));
 sky130_fd_sc_hd__a22o_1 _4380_ (.A1(\BitStream_buffer.BS_buffer[39] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[40] ),
    .X(_1165_));
 sky130_fd_sc_hd__or4_1 _4381_ (.A(_1162_),
    .B(_1163_),
    .C(_1164_),
    .D(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__o22ai_1 _4382_ (.A1(_0499_),
    .A2(_2941_),
    .B1(_2963_),
    .B2(_2945_),
    .Y(_1167_));
 sky130_fd_sc_hd__a221oi_1 _4383_ (.A1(\BitStream_buffer.BS_buffer[51] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[52] ),
    .B2(_2938_),
    .C1(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__o22ai_1 _4384_ (.A1(_2975_),
    .A2(_2955_),
    .B1(_0619_),
    .B2(_2959_),
    .Y(_1169_));
 sky130_fd_sc_hd__a221oi_1 _4385_ (.A1(\BitStream_buffer.BS_buffer[47] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[48] ),
    .B2(_2952_),
    .C1(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__nand3b_1 _4386_ (.A_N(_1166_),
    .B(_1168_),
    .C(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__o22ai_1 _4387_ (.A1(_0505_),
    .A2(_2967_),
    .B1(_2996_),
    .B2(_2970_),
    .Y(_1172_));
 sky130_fd_sc_hd__o22ai_1 _4388_ (.A1(_2999_),
    .A2(_2974_),
    .B1(_0858_),
    .B2(_2977_),
    .Y(_1173_));
 sky130_fd_sc_hd__a22o_1 _4389_ (.A1(\BitStream_buffer.BS_buffer[61] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[62] ),
    .X(_1174_));
 sky130_fd_sc_hd__a22o_1 _4390_ (.A1(\BitStream_buffer.BS_buffer[55] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[56] ),
    .X(_1175_));
 sky130_fd_sc_hd__or4_1 _4391_ (.A(_1172_),
    .B(_1173_),
    .C(_1174_),
    .D(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__o22ai_1 _4392_ (.A1(_0411_),
    .A2(_2998_),
    .B1(_2652_),
    .B2(_3001_),
    .Y(_1177_));
 sky130_fd_sc_hd__a221oi_1 _4393_ (.A1(\BitStream_buffer.BS_buffer[63] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[64] ),
    .B2(_2995_),
    .C1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__a2bb2o_1 _4394_ (.A1_N(_2664_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[70] ),
    .B2(_3014_),
    .X(_1179_));
 sky130_fd_sc_hd__a221oi_1 _4395_ (.A1(\BitStream_buffer.BS_buffer[67] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[68] ),
    .B2(_3008_),
    .C1(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__nand3b_1 _4396_ (.A_N(_1176_),
    .B(_1178_),
    .C(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__nor2_1 _4397_ (.A(_0514_),
    .B(_3022_),
    .Y(_1182_));
 sky130_fd_sc_hd__o22ai_1 _4398_ (.A1(_3056_),
    .A2(_3026_),
    .B1(_0648_),
    .B2(_3030_),
    .Y(_1183_));
 sky130_fd_sc_hd__a22o_1 _4399_ (.A1(_0650_),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_0770_),
    .X(_1184_));
 sky130_fd_sc_hd__a22o_1 _4400_ (.A1(_0325_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_0527_),
    .X(_1185_));
 sky130_fd_sc_hd__or4_1 _4401_ (.A(_1182_),
    .B(_1183_),
    .C(_1184_),
    .D(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__a22o_1 _4402_ (.A1(\BitStream_buffer.BS_buffer[19] ),
    .A2(_3048_),
    .B1(_3050_),
    .B2(\BitStream_buffer.BS_buffer[20] ),
    .X(_1187_));
 sky130_fd_sc_hd__o22ai_1 _4403_ (.A1(_0358_),
    .A2(_3055_),
    .B1(_0660_),
    .B2(_3058_),
    .Y(_1188_));
 sky130_fd_sc_hd__o22ai_1 _4404_ (.A1(_0373_),
    .A2(_3062_),
    .B1(_0646_),
    .B2(_0323_),
    .Y(_1189_));
 sky130_fd_sc_hd__a22o_1 _4405_ (.A1(_0363_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(\BitStream_buffer.BS_buffer[15] ),
    .X(_1190_));
 sky130_fd_sc_hd__or4_1 _4406_ (.A(_1187_),
    .B(_1188_),
    .C(_1189_),
    .D(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__nor2_1 _4407_ (.A(_1186_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__o22ai_1 _4408_ (.A1(_2917_),
    .A2(_0344_),
    .B1(_0663_),
    .B2(_0347_),
    .Y(_1193_));
 sky130_fd_sc_hd__a221oi_1 _4409_ (.A1(\BitStream_buffer.BS_buffer[32] ),
    .A2(_0340_),
    .B1(\BitStream_buffer.BS_buffer[31] ),
    .B2(_0337_),
    .C1(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__o22ai_1 _4410_ (.A1(_0388_),
    .A2(_0357_),
    .B1(_0654_),
    .B2(_0360_),
    .Y(_1195_));
 sky130_fd_sc_hd__a221oi_1 _4411_ (.A1(\BitStream_buffer.BS_buffer[27] ),
    .A2(_0351_),
    .B1(\BitStream_buffer.BS_buffer[28] ),
    .B2(_0354_),
    .C1(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__o22ai_1 _4412_ (.A1(_0345_),
    .A2(_0372_),
    .B1(_0657_),
    .B2(_0375_),
    .Y(_1197_));
 sky130_fd_sc_hd__a221oi_1 _4413_ (.A1(\BitStream_buffer.BS_buffer[23] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[24] ),
    .B2(_0369_),
    .C1(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__o22ai_1 _4414_ (.A1(_0486_),
    .A2(_0386_),
    .B1(_2905_),
    .B2(_0390_),
    .Y(_1199_));
 sky130_fd_sc_hd__a221oi_1 _4415_ (.A1(\BitStream_buffer.BS_buffer[35] ),
    .A2(_0379_),
    .B1(\BitStream_buffer.BS_buffer[36] ),
    .B2(_0383_),
    .C1(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__and4_1 _4416_ (.A(_1194_),
    .B(_1196_),
    .C(_1198_),
    .D(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__nand2_1 _4417_ (.A(_1192_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__nor3_1 _4418_ (.A(_1171_),
    .B(_1181_),
    .C(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_0399_),
    .B(\BitStream_buffer.BS_buffer[7] ),
    .Y(_1204_));
 sky130_fd_sc_hd__nand3_1 _4420_ (.A(_1161_),
    .B(_1203_),
    .C(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__inv_2 _4421_ (.A(\BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_1206_));
 sky130_fd_sc_hd__a21oi_1 _4422_ (.A1(_1206_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1207_));
 sky130_fd_sc_hd__o21a_1 _4423_ (.A1(_2599_),
    .A2(_1205_),
    .B1(_1207_),
    .X(_0314_));
 sky130_fd_sc_hd__o22ai_1 _4424_ (.A1(_2742_),
    .A2(_2630_),
    .B1(_0686_),
    .B2(_2637_),
    .Y(_1208_));
 sky130_fd_sc_hd__a221oi_1 _4425_ (.A1(\BitStream_buffer.BS_buffer[82] ),
    .A2(_2617_),
    .B1(\BitStream_buffer.BS_buffer[83] ),
    .B2(_2624_),
    .C1(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2_1 _4426_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[74] ),
    .Y(_1210_));
 sky130_fd_sc_hd__or2_1 _4427_ (.A(_2625_),
    .B(_2656_),
    .X(_1211_));
 sky130_fd_sc_hd__or2_1 _4428_ (.A(_0549_),
    .B(_2661_),
    .X(_1212_));
 sky130_fd_sc_hd__o2111a_1 _4429_ (.A1(_2631_),
    .A2(_2646_),
    .B1(_1210_),
    .C1(_1211_),
    .D1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__o22ai_1 _4430_ (.A1(_2694_),
    .A2(_2670_),
    .B1(_2698_),
    .B2(_2675_),
    .Y(_1214_));
 sky130_fd_sc_hd__a22o_1 _4431_ (.A1(\BitStream_buffer.BS_buffer[78] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[79] ),
    .X(_1215_));
 sky130_fd_sc_hd__nor2_1 _4432_ (.A(_1214_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__o22ai_1 _4433_ (.A1(_2769_),
    .A2(_2697_),
    .B1(_0434_),
    .B2(_2702_),
    .Y(_1217_));
 sky130_fd_sc_hd__a221oi_1 _4434_ (.A1(_2762_),
    .A2(_2689_),
    .B1(_2756_),
    .B2(_2693_),
    .C1(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__and4_1 _4435_ (.A(_1209_),
    .B(_1213_),
    .C(_1216_),
    .D(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__or2_1 _4436_ (.A(_2795_),
    .B(_2717_),
    .X(_1220_));
 sky130_fd_sc_hd__nand2_1 _4437_ (.A(_2720_),
    .B(_2804_),
    .Y(_1221_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(_2724_),
    .B(_2800_),
    .Y(_1222_));
 sky130_fd_sc_hd__o2111a_1 _4439_ (.A1(_2806_),
    .A2(_2713_),
    .B1(_1220_),
    .C1(_1221_),
    .D1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__o22ai_1 _4440_ (.A1(_2822_),
    .A2(_2735_),
    .B1(_0450_),
    .B2(_2739_),
    .Y(_1224_));
 sky130_fd_sc_hd__a221oi_1 _4441_ (.A1(_2816_),
    .A2(_2729_),
    .B1(\BitStream_buffer.BS_buffer[103] ),
    .B2(_2732_),
    .C1(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(_2746_),
    .B(_2721_),
    .Y(_1226_));
 sky130_fd_sc_hd__nand2_1 _4443_ (.A(_2749_),
    .B(_2725_),
    .Y(_1227_));
 sky130_fd_sc_hd__or2_1 _4444_ (.A(_2715_),
    .B(_2753_),
    .X(_1228_));
 sky130_fd_sc_hd__o2111a_1 _4445_ (.A1(_2707_),
    .A2(_2744_),
    .B1(_1226_),
    .C1(_1227_),
    .D1(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__nand2_1 _4446_ (.A(_2761_),
    .B(\BitStream_buffer.BS_buffer[94] ),
    .Y(_1230_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(_2765_),
    .B(_2736_),
    .Y(_1231_));
 sky130_fd_sc_hd__or2_1 _4448_ (.A(_2733_),
    .B(_2771_),
    .X(_1232_));
 sky130_fd_sc_hd__o2111a_1 _4449_ (.A1(_0568_),
    .A2(_2759_),
    .B1(_1230_),
    .C1(_1231_),
    .D1(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__and4_1 _4450_ (.A(_1223_),
    .B(_1225_),
    .C(_1229_),
    .D(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__or2_1 _4451_ (.A(_2894_),
    .B(_2784_),
    .X(_1235_));
 sky130_fd_sc_hd__nand2_1 _4452_ (.A(_2787_),
    .B(\BitStream_buffer.BS_buffer[114] ),
    .Y(_1236_));
 sky130_fd_sc_hd__nand2_1 _4453_ (.A(_2791_),
    .B(\BitStream_buffer.BS_buffer[112] ),
    .Y(_1237_));
 sky130_fd_sc_hd__o2111a_1 _4454_ (.A1(_2898_),
    .A2(_2780_),
    .B1(_1235_),
    .C1(_1236_),
    .D1(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__nand2_1 _4455_ (.A(_2799_),
    .B(_2792_),
    .Y(_1239_));
 sky130_fd_sc_hd__nand2_1 _4456_ (.A(_2803_),
    .B(_2788_),
    .Y(_1240_));
 sky130_fd_sc_hd__or2_1 _4457_ (.A(_2775_),
    .B(_2808_),
    .X(_1241_));
 sky130_fd_sc_hd__o2111a_1 _4458_ (.A1(_2782_),
    .A2(_2797_),
    .B1(_1239_),
    .C1(_1240_),
    .D1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__nand2_1 _4459_ (.A(_2815_),
    .B(_2836_),
    .Y(_1243_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_2819_),
    .B(_2832_),
    .Y(_1244_));
 sky130_fd_sc_hd__or2_1 _4461_ (.A(_2839_),
    .B(_2824_),
    .X(_1245_));
 sky130_fd_sc_hd__o2111a_1 _4462_ (.A1(_2827_),
    .A2(_2813_),
    .B1(_1243_),
    .C1(_1244_),
    .D1(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__nand2_1 _4463_ (.A(_2831_),
    .B(\BitStream_buffer.BS_buffer[116] ),
    .Y(_1247_));
 sky130_fd_sc_hd__nand2_1 _4464_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[118] ),
    .Y(_1248_));
 sky130_fd_sc_hd__or2_1 _4465_ (.A(_2867_),
    .B(_2841_),
    .X(_1249_));
 sky130_fd_sc_hd__o2111a_1 _4466_ (.A1(_0601_),
    .A2(_2829_),
    .B1(_1247_),
    .C1(_1248_),
    .D1(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__and4_1 _4467_ (.A(_1238_),
    .B(_1242_),
    .C(_1246_),
    .D(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__or2_1 _4468_ (.A(_3018_),
    .B(_2852_),
    .X(_1252_));
 sky130_fd_sc_hd__nand2_1 _4469_ (.A(_2856_),
    .B(_3039_),
    .Y(_1253_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_2859_),
    .B(_0400_),
    .Y(_1254_));
 sky130_fd_sc_hd__o2111a_1 _4471_ (.A1(_0638_),
    .A2(_2849_),
    .B1(_1252_),
    .C1(_1253_),
    .D1(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__o22ai_1 _4472_ (.A1(_2880_),
    .A2(_2869_),
    .B1(_2883_),
    .B2(_2872_),
    .Y(_1256_));
 sky130_fd_sc_hd__a221oi_1 _4473_ (.A1(\BitStream_buffer.BS_buffer[126] ),
    .A2(_2863_),
    .B1(\BitStream_buffer.BS_buffer[127] ),
    .B2(_2866_),
    .C1(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__o22ai_1 _4474_ (.A1(_0869_),
    .A2(_2882_),
    .B1(_0761_),
    .B2(_2885_),
    .Y(_1258_));
 sky130_fd_sc_hd__a221oi_1 _4475_ (.A1(_0516_),
    .A2(_2876_),
    .B1(\BitStream_buffer.BS_buffer[7] ),
    .B2(_2879_),
    .C1(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_1 _4476_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[122] ),
    .Y(_1260_));
 sky130_fd_sc_hd__or2_1 _4477_ (.A(_2845_),
    .B(_2896_),
    .X(_1261_));
 sky130_fd_sc_hd__or2_1 _4478_ (.A(_2850_),
    .B(_2900_),
    .X(_1262_));
 sky130_fd_sc_hd__o2111a_1 _4479_ (.A1(_0727_),
    .A2(_2890_),
    .B1(_1260_),
    .C1(_1261_),
    .D1(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__and4_1 _4480_ (.A(_1255_),
    .B(_1257_),
    .C(_1259_),
    .D(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__and4_1 _4481_ (.A(_1219_),
    .B(_1234_),
    .C(_1251_),
    .D(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__o22ai_1 _4482_ (.A1(_0622_),
    .A2(_2909_),
    .B1(_0495_),
    .B2(_2912_),
    .Y(_1266_));
 sky130_fd_sc_hd__o22ai_1 _4483_ (.A1(_2953_),
    .A2(_2916_),
    .B1(_2956_),
    .B2(_2920_),
    .Y(_1267_));
 sky130_fd_sc_hd__a22o_1 _4484_ (.A1(\BitStream_buffer.BS_buffer[46] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[47] ),
    .X(_1268_));
 sky130_fd_sc_hd__a22o_1 _4485_ (.A1(\BitStream_buffer.BS_buffer[40] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[41] ),
    .X(_1269_));
 sky130_fd_sc_hd__or4_1 _4486_ (.A(_1266_),
    .B(_1267_),
    .C(_1268_),
    .D(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__o22ai_1 _4487_ (.A1(_0626_),
    .A2(_2941_),
    .B1(_0499_),
    .B2(_2945_),
    .Y(_1271_));
 sky130_fd_sc_hd__a221oi_2 _4488_ (.A1(\BitStream_buffer.BS_buffer[52] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[53] ),
    .B2(_2938_),
    .C1(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__o22ai_1 _4489_ (.A1(_2972_),
    .A2(_2955_),
    .B1(_2975_),
    .B2(_2959_),
    .Y(_1273_));
 sky130_fd_sc_hd__a221oi_1 _4490_ (.A1(\BitStream_buffer.BS_buffer[48] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[49] ),
    .B2(_2952_),
    .C1(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__nand3b_1 _4491_ (.A_N(_1270_),
    .B(_1272_),
    .C(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__o22ai_1 _4492_ (.A1(_0632_),
    .A2(_2967_),
    .B1(_0505_),
    .B2(_2970_),
    .Y(_1276_));
 sky130_fd_sc_hd__o22ai_1 _4493_ (.A1(_2996_),
    .A2(_2974_),
    .B1(_2999_),
    .B2(_2977_),
    .Y(_1277_));
 sky130_fd_sc_hd__a22o_1 _4494_ (.A1(\BitStream_buffer.BS_buffer[62] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[63] ),
    .X(_1278_));
 sky130_fd_sc_hd__a22o_1 _4495_ (.A1(\BitStream_buffer.BS_buffer[56] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[57] ),
    .X(_1279_));
 sky130_fd_sc_hd__or4_1 _4496_ (.A(_1276_),
    .B(_1277_),
    .C(_1278_),
    .D(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__o22ai_1 _4497_ (.A1(_2658_),
    .A2(_2998_),
    .B1(_0411_),
    .B2(_3001_),
    .Y(_1281_));
 sky130_fd_sc_hd__a221oi_1 _4498_ (.A1(\BitStream_buffer.BS_buffer[64] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[65] ),
    .B2(_2995_),
    .C1(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__a2bb2o_1 _4499_ (.A1_N(_0415_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[71] ),
    .B2(_3014_),
    .X(_1283_));
 sky130_fd_sc_hd__a221oi_1 _4500_ (.A1(\BitStream_buffer.BS_buffer[68] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[69] ),
    .B2(_3008_),
    .C1(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__nand3b_1 _4501_ (.A_N(_1280_),
    .B(_1282_),
    .C(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__nor2_1 _4502_ (.A(_0640_),
    .B(_3022_),
    .Y(_1286_));
 sky130_fd_sc_hd__o22ai_1 _4503_ (.A1(_3053_),
    .A2(_3026_),
    .B1(_3056_),
    .B2(_3030_),
    .Y(_1287_));
 sky130_fd_sc_hd__a22o_1 _4504_ (.A1(_0770_),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_3051_),
    .X(_1288_));
 sky130_fd_sc_hd__a22o_1 _4505_ (.A1(_0527_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_0650_),
    .X(_1289_));
 sky130_fd_sc_hd__or4_1 _4506_ (.A(_1286_),
    .B(_1287_),
    .C(_1288_),
    .D(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__a22o_1 _4507_ (.A1(\BitStream_buffer.BS_buffer[20] ),
    .A2(_3048_),
    .B1(_3050_),
    .B2(\BitStream_buffer.BS_buffer[21] ),
    .X(_1291_));
 sky130_fd_sc_hd__o22ai_1 _4508_ (.A1(_0355_),
    .A2(_3055_),
    .B1(_0358_),
    .B2(_3058_),
    .Y(_1292_));
 sky130_fd_sc_hd__o22ai_1 _4509_ (.A1(_0370_),
    .A2(_3062_),
    .B1(_0373_),
    .B2(_0323_),
    .Y(_1293_));
 sky130_fd_sc_hd__a22o_1 _4510_ (.A1(_0366_),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0363_),
    .X(_1294_));
 sky130_fd_sc_hd__or4_1 _4511_ (.A(_1291_),
    .B(_1292_),
    .C(_1293_),
    .D(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__nor2_1 _4512_ (.A(_1290_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__o22ai_1 _4513_ (.A1(_2914_),
    .A2(_0344_),
    .B1(_2917_),
    .B2(_0347_),
    .Y(_1297_));
 sky130_fd_sc_hd__a221oi_1 _4514_ (.A1(\BitStream_buffer.BS_buffer[32] ),
    .A2(_0337_),
    .B1(\BitStream_buffer.BS_buffer[33] ),
    .B2(_0341_),
    .C1(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__o22ai_1 _4515_ (.A1(_0384_),
    .A2(_0357_),
    .B1(_0388_),
    .B2(_0360_),
    .Y(_1299_));
 sky130_fd_sc_hd__a221oi_1 _4516_ (.A1(\BitStream_buffer.BS_buffer[28] ),
    .A2(_0351_),
    .B1(_0380_),
    .B2(_0354_),
    .C1(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__o22ai_1 _4517_ (.A1(_0342_),
    .A2(_0372_),
    .B1(_0345_),
    .B2(_0375_),
    .Y(_1301_));
 sky130_fd_sc_hd__a221oi_1 _4518_ (.A1(\BitStream_buffer.BS_buffer[24] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[25] ),
    .B2(_0369_),
    .C1(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__o22ai_1 _4519_ (.A1(_0613_),
    .A2(_0386_),
    .B1(_0486_),
    .B2(_0390_),
    .Y(_1303_));
 sky130_fd_sc_hd__a221oi_1 _4520_ (.A1(\BitStream_buffer.BS_buffer[36] ),
    .A2(_0379_),
    .B1(\BitStream_buffer.BS_buffer[37] ),
    .B2(_0383_),
    .C1(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__and4_1 _4521_ (.A(_1298_),
    .B(_1300_),
    .C(_1302_),
    .D(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__nand2_1 _4522_ (.A(_1296_),
    .B(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__nor3_1 _4523_ (.A(_1275_),
    .B(_1285_),
    .C(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_0399_),
    .B(_0330_),
    .Y(_1308_));
 sky130_fd_sc_hd__nand3_1 _4525_ (.A(_1265_),
    .B(_1307_),
    .C(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__inv_2 _4526_ (.A(\BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_1310_));
 sky130_fd_sc_hd__a21oi_1 _4527_ (.A1(_1310_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1311_));
 sky130_fd_sc_hd__o21a_1 _4528_ (.A1(_2599_),
    .A2(_1309_),
    .B1(_1311_),
    .X(_0313_));
 sky130_fd_sc_hd__o22ai_1 _4529_ (.A1(_0431_),
    .A2(_2630_),
    .B1(_2742_),
    .B2(_2637_),
    .Y(_1312_));
 sky130_fd_sc_hd__a221oi_1 _4530_ (.A1(\BitStream_buffer.BS_buffer[83] ),
    .A2(_2617_),
    .B1(_2766_),
    .B2(_2624_),
    .C1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2_1 _4531_ (.A(_2650_),
    .B(\BitStream_buffer.BS_buffer[75] ),
    .Y(_1314_));
 sky130_fd_sc_hd__or2_1 _4532_ (.A(_0407_),
    .B(_2656_),
    .X(_1315_));
 sky130_fd_sc_hd__or2_1 _4533_ (.A(_2698_),
    .B(_2661_),
    .X(_1316_));
 sky130_fd_sc_hd__o2111a_1 _4534_ (.A1(_2625_),
    .A2(_2646_),
    .B1(_1314_),
    .C1(_1315_),
    .D1(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__o22ai_1 _4535_ (.A1(_0419_),
    .A2(_2670_),
    .B1(_2694_),
    .B2(_2675_),
    .Y(_1318_));
 sky130_fd_sc_hd__a22o_1 _4536_ (.A1(\BitStream_buffer.BS_buffer[79] ),
    .A2(_2679_),
    .B1(_2682_),
    .B2(\BitStream_buffer.BS_buffer[80] ),
    .X(_1319_));
 sky130_fd_sc_hd__nor2_1 _4537_ (.A(_1318_),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__o22ai_1 _4538_ (.A1(_0440_),
    .A2(_2697_),
    .B1(_2769_),
    .B2(_2702_),
    .Y(_1321_));
 sky130_fd_sc_hd__a221oi_1 _4539_ (.A1(_2756_),
    .A2(_2689_),
    .B1(_2725_),
    .B2(_2693_),
    .C1(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__and4_1 _4540_ (.A(_1313_),
    .B(_1317_),
    .C(_1320_),
    .D(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__or2_1 _4541_ (.A(_0450_),
    .B(_2717_),
    .X(_1324_));
 sky130_fd_sc_hd__nand2_1 _4542_ (.A(_2720_),
    .B(\BitStream_buffer.BS_buffer[99] ),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _4543_ (.A(_2724_),
    .B(\BitStream_buffer.BS_buffer[97] ),
    .Y(_1326_));
 sky130_fd_sc_hd__o2111a_1 _4544_ (.A1(_0453_),
    .A2(_2713_),
    .B1(_1324_),
    .C1(_1325_),
    .D1(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__o22ai_1 _4545_ (.A1(_0459_),
    .A2(_2735_),
    .B1(_2822_),
    .B2(_2739_),
    .Y(_1328_));
 sky130_fd_sc_hd__a221oi_1 _4546_ (.A1(\BitStream_buffer.BS_buffer[103] ),
    .A2(_2729_),
    .B1(_2792_),
    .B2(_2732_),
    .C1(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__nand2_1 _4547_ (.A(_2746_),
    .B(_2714_),
    .Y(_1330_));
 sky130_fd_sc_hd__nand2_1 _4548_ (.A(_2749_),
    .B(_2706_),
    .Y(_1331_));
 sky130_fd_sc_hd__or2_1 _4549_ (.A(_2737_),
    .B(_2753_),
    .X(_1332_));
 sky130_fd_sc_hd__o2111a_1 _4550_ (.A1(_0423_),
    .A2(_2744_),
    .B1(_1330_),
    .C1(_1331_),
    .D1(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__nand2_1 _4551_ (.A(_2761_),
    .B(\BitStream_buffer.BS_buffer[95] ),
    .Y(_1334_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(_2765_),
    .B(\BitStream_buffer.BS_buffer[93] ),
    .Y(_1335_));
 sky130_fd_sc_hd__or2_1 _4553_ (.A(_0428_),
    .B(_2771_),
    .X(_1336_));
 sky130_fd_sc_hd__o2111a_1 _4554_ (.A1(_0694_),
    .A2(_2759_),
    .B1(_1334_),
    .C1(_1335_),
    .D1(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__and4_1 _4555_ (.A(_1327_),
    .B(_1329_),
    .C(_1333_),
    .D(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__or2_1 _4556_ (.A(_2870_),
    .B(_2784_),
    .X(_1339_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_2787_),
    .B(\BitStream_buffer.BS_buffer[115] ),
    .Y(_1340_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_2791_),
    .B(\BitStream_buffer.BS_buffer[113] ),
    .Y(_1341_));
 sky130_fd_sc_hd__o2111a_1 _4559_ (.A1(_0481_),
    .A2(_2780_),
    .B1(_1339_),
    .C1(_1340_),
    .D1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_2799_),
    .B(\BitStream_buffer.BS_buffer[105] ),
    .Y(_1343_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_2803_),
    .B(_2781_),
    .Y(_1344_));
 sky130_fd_sc_hd__or2_1 _4562_ (.A(_0444_),
    .B(_2808_),
    .X(_1345_));
 sky130_fd_sc_hd__o2111a_1 _4563_ (.A1(_0445_),
    .A2(_2797_),
    .B1(_1343_),
    .C1(_1344_),
    .D1(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_2815_),
    .B(\BitStream_buffer.BS_buffer[111] ),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2_1 _4565_ (.A(_2819_),
    .B(_2838_),
    .Y(_1348_));
 sky130_fd_sc_hd__or2_1 _4566_ (.A(_0464_),
    .B(_2824_),
    .X(_1349_));
 sky130_fd_sc_hd__o2111a_1 _4567_ (.A1(_2888_),
    .A2(_2813_),
    .B1(_1347_),
    .C1(_1348_),
    .D1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__nand2_1 _4568_ (.A(_2831_),
    .B(\BitStream_buffer.BS_buffer[117] ),
    .Y(_1351_));
 sky130_fd_sc_hd__nand2_1 _4569_ (.A(_2835_),
    .B(\BitStream_buffer.BS_buffer[119] ),
    .Y(_1352_));
 sky130_fd_sc_hd__or2_1 _4570_ (.A(_0473_),
    .B(_2841_),
    .X(_1353_));
 sky130_fd_sc_hd__o2111a_1 _4571_ (.A1(_0727_),
    .A2(_2829_),
    .B1(_1351_),
    .C1(_1352_),
    .D1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__and4_1 _4572_ (.A(_1342_),
    .B(_1346_),
    .C(_1350_),
    .D(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__or2_1 _4573_ (.A(_0512_),
    .B(_2852_),
    .X(_1356_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(_2856_),
    .B(_3044_),
    .Y(_1357_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_2859_),
    .B(\BitStream_buffer.BS_buffer[1] ),
    .Y(_1358_));
 sky130_fd_sc_hd__o2111a_1 _4576_ (.A1(_0761_),
    .A2(_2849_),
    .B1(_1356_),
    .C1(_1357_),
    .D1(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__o22ai_1 _4577_ (.A1(_0476_),
    .A2(_2869_),
    .B1(_2880_),
    .B2(_2872_),
    .Y(_1360_));
 sky130_fd_sc_hd__a221oi_1 _4578_ (.A1(_0400_),
    .A2(_2865_),
    .B1(\BitStream_buffer.BS_buffer[127] ),
    .B2(_2863_),
    .C1(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__o22ai_1 _4579_ (.A1(_3027_),
    .A2(_2882_),
    .B1(_0869_),
    .B2(_2885_),
    .Y(_1362_));
 sky130_fd_sc_hd__a221oi_1 _4580_ (.A1(\BitStream_buffer.BS_buffer[7] ),
    .A2(_2876_),
    .B1(_0330_),
    .B2(_2879_),
    .C1(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(_2892_),
    .B(\BitStream_buffer.BS_buffer[123] ),
    .Y(_1364_));
 sky130_fd_sc_hd__or2_1 _4582_ (.A(_2883_),
    .B(_2896_),
    .X(_1365_));
 sky130_fd_sc_hd__or2_1 _4583_ (.A(_0468_),
    .B(_2900_),
    .X(_1366_));
 sky130_fd_sc_hd__o2111a_1 _4584_ (.A1(_2850_),
    .A2(_2890_),
    .B1(_1364_),
    .C1(_1365_),
    .D1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__and4_1 _4585_ (.A(_1359_),
    .B(_1361_),
    .C(_1363_),
    .D(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__and4_1 _4586_ (.A(_1323_),
    .B(_1338_),
    .C(_1355_),
    .D(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__o22ai_1 _4587_ (.A1(_2942_),
    .A2(_2909_),
    .B1(_0622_),
    .B2(_2912_),
    .Y(_1370_));
 sky130_fd_sc_hd__o22ai_1 _4588_ (.A1(_0495_),
    .A2(_2916_),
    .B1(_2953_),
    .B2(_2920_),
    .Y(_1371_));
 sky130_fd_sc_hd__a22o_1 _4589_ (.A1(\BitStream_buffer.BS_buffer[47] ),
    .A2(_2924_),
    .B1(_2926_),
    .B2(\BitStream_buffer.BS_buffer[48] ),
    .X(_1372_));
 sky130_fd_sc_hd__a22o_1 _4590_ (.A1(\BitStream_buffer.BS_buffer[41] ),
    .A2(_2929_),
    .B1(_2931_),
    .B2(\BitStream_buffer.BS_buffer[42] ),
    .X(_1373_));
 sky130_fd_sc_hd__or4_1 _4591_ (.A(_1370_),
    .B(_1371_),
    .C(_1372_),
    .D(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__o22ai_1 _4592_ (.A1(_0750_),
    .A2(_2941_),
    .B1(_0626_),
    .B2(_2945_),
    .Y(_1375_));
 sky130_fd_sc_hd__a221oi_1 _4593_ (.A1(\BitStream_buffer.BS_buffer[53] ),
    .A2(_2935_),
    .B1(\BitStream_buffer.BS_buffer[54] ),
    .B2(_2938_),
    .C1(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__o22ai_1 _4594_ (.A1(_2968_),
    .A2(_2955_),
    .B1(_2972_),
    .B2(_2959_),
    .Y(_1377_));
 sky130_fd_sc_hd__a221oi_1 _4595_ (.A1(\BitStream_buffer.BS_buffer[49] ),
    .A2(_2949_),
    .B1(\BitStream_buffer.BS_buffer[50] ),
    .B2(_2952_),
    .C1(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand3b_1 _4596_ (.A_N(_1374_),
    .B(_1376_),
    .C(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__o22ai_1 _4597_ (.A1(_3009_),
    .A2(_2967_),
    .B1(_0632_),
    .B2(_2970_),
    .Y(_1380_));
 sky130_fd_sc_hd__o22ai_1 _4598_ (.A1(_0505_),
    .A2(_2974_),
    .B1(_2996_),
    .B2(_2977_),
    .Y(_1381_));
 sky130_fd_sc_hd__a22o_1 _4599_ (.A1(\BitStream_buffer.BS_buffer[63] ),
    .A2(_2981_),
    .B1(_2983_),
    .B2(\BitStream_buffer.BS_buffer[64] ),
    .X(_1382_));
 sky130_fd_sc_hd__a22o_1 _4600_ (.A1(\BitStream_buffer.BS_buffer[57] ),
    .A2(_2986_),
    .B1(_2988_),
    .B2(\BitStream_buffer.BS_buffer[58] ),
    .X(_1383_));
 sky130_fd_sc_hd__or4_1 _4601_ (.A(_1380_),
    .B(_1381_),
    .C(_1382_),
    .D(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__o22ai_1 _4602_ (.A1(_2671_),
    .A2(_2998_),
    .B1(_2658_),
    .B2(_3001_),
    .Y(_1385_));
 sky130_fd_sc_hd__a221oi_1 _4603_ (.A1(\BitStream_buffer.BS_buffer[65] ),
    .A2(_2992_),
    .B1(\BitStream_buffer.BS_buffer[66] ),
    .B2(_2995_),
    .C1(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__a2bb2o_1 _4604_ (.A1_N(_0556_),
    .A2_N(_3011_),
    .B1(\BitStream_buffer.BS_buffer[72] ),
    .B2(_3014_),
    .X(_1387_));
 sky130_fd_sc_hd__a221oi_1 _4605_ (.A1(\BitStream_buffer.BS_buffer[69] ),
    .A2(_3005_),
    .B1(\BitStream_buffer.BS_buffer[70] ),
    .B2(_3008_),
    .C1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__nand3b_1 _4606_ (.A_N(_1384_),
    .B(_1386_),
    .C(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__nor2_1 _4607_ (.A(_3063_),
    .B(_3022_),
    .Y(_1390_));
 sky130_fd_sc_hd__o22ai_1 _4608_ (.A1(_0523_),
    .A2(_3026_),
    .B1(_3053_),
    .B2(_3030_),
    .Y(_1391_));
 sky130_fd_sc_hd__a22o_1 _4609_ (.A1(_3051_),
    .A2(_3034_),
    .B1(_3036_),
    .B2(_0521_),
    .X(_1392_));
 sky130_fd_sc_hd__a22o_1 _4610_ (.A1(_0650_),
    .A2(_3041_),
    .B1(_3043_),
    .B2(_0770_),
    .X(_1393_));
 sky130_fd_sc_hd__or4_1 _4611_ (.A(_1390_),
    .B(_1391_),
    .C(_1392_),
    .D(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__a22o_1 _4612_ (.A1(\BitStream_buffer.BS_buffer[21] ),
    .A2(_3048_),
    .B1(_3050_),
    .B2(\BitStream_buffer.BS_buffer[22] ),
    .X(_1395_));
 sky130_fd_sc_hd__o22ai_1 _4613_ (.A1(_0534_),
    .A2(_3055_),
    .B1(_0355_),
    .B2(_3058_),
    .Y(_1396_));
 sky130_fd_sc_hd__o22ai_1 _4614_ (.A1(_0537_),
    .A2(_3062_),
    .B1(_0370_),
    .B2(_0323_),
    .Y(_1397_));
 sky130_fd_sc_hd__a22o_1 _4615_ (.A1(\BitStream_buffer.BS_buffer[18] ),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0366_),
    .X(_1398_));
 sky130_fd_sc_hd__or4_1 _4616_ (.A(_1395_),
    .B(_1396_),
    .C(_1397_),
    .D(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__nor2_1 _4617_ (.A(_1394_),
    .B(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__o22ai_1 _4618_ (.A1(_2910_),
    .A2(_0344_),
    .B1(_2914_),
    .B2(_0347_),
    .Y(_1401_));
 sky130_fd_sc_hd__a221oi_1 _4619_ (.A1(\BitStream_buffer.BS_buffer[33] ),
    .A2(_0337_),
    .B1(\BitStream_buffer.BS_buffer[34] ),
    .B2(_0341_),
    .C1(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__o22ai_1 _4620_ (.A1(_0540_),
    .A2(_0357_),
    .B1(_0384_),
    .B2(_0360_),
    .Y(_1403_));
 sky130_fd_sc_hd__a221oi_1 _4621_ (.A1(_0380_),
    .A2(_0350_),
    .B1(_0387_),
    .B2(_0354_),
    .C1(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__o22ai_1 _4622_ (.A1(_0531_),
    .A2(_0372_),
    .B1(_0342_),
    .B2(_0375_),
    .Y(_1405_));
 sky130_fd_sc_hd__a221oi_1 _4623_ (.A1(\BitStream_buffer.BS_buffer[25] ),
    .A2(_0365_),
    .B1(\BitStream_buffer.BS_buffer[26] ),
    .B2(_0369_),
    .C1(_1405_),
    .Y(_1406_));
 sky130_fd_sc_hd__o22ai_1 _4624_ (.A1(_0739_),
    .A2(_0386_),
    .B1(_0613_),
    .B2(_0390_),
    .Y(_1407_));
 sky130_fd_sc_hd__a221oi_1 _4625_ (.A1(\BitStream_buffer.BS_buffer[37] ),
    .A2(_0379_),
    .B1(\BitStream_buffer.BS_buffer[38] ),
    .B2(_0383_),
    .C1(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__and4_1 _4626_ (.A(_1402_),
    .B(_1404_),
    .C(_1406_),
    .D(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__nand2_1 _4627_ (.A(_1400_),
    .B(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__nor3_1 _4628_ (.A(_1379_),
    .B(_1389_),
    .C(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(_0399_),
    .B(_0325_),
    .Y(_1412_));
 sky130_fd_sc_hd__nand3_1 _4630_ (.A(_1369_),
    .B(_1411_),
    .C(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__inv_2 _4631_ (.A(\BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_1414_));
 sky130_fd_sc_hd__a21oi_1 _4632_ (.A1(_1414_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1415_));
 sky130_fd_sc_hd__o21a_1 _4633_ (.A1(_2599_),
    .A2(_1413_),
    .B1(_1415_),
    .X(_0312_));
 sky130_fd_sc_hd__o22ai_1 _4634_ (.A1(_2751_),
    .A2(_2629_),
    .B1(_0431_),
    .B2(_2636_),
    .Y(_1416_));
 sky130_fd_sc_hd__a221oi_1 _4635_ (.A1(_2766_),
    .A2(_2616_),
    .B1(_2768_),
    .B2(_2623_),
    .C1(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _4636_ (.A(_2649_),
    .B(\BitStream_buffer.BS_buffer[76] ),
    .Y(_1418_));
 sky130_fd_sc_hd__or2_1 _4637_ (.A(_0549_),
    .B(_2655_),
    .X(_1419_));
 sky130_fd_sc_hd__or2_1 _4638_ (.A(_2694_),
    .B(_2660_),
    .X(_1420_));
 sky130_fd_sc_hd__o2111a_1 _4639_ (.A1(_0407_),
    .A2(_2645_),
    .B1(_1418_),
    .C1(_1419_),
    .D1(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__o22ai_1 _4640_ (.A1(_0560_),
    .A2(_2669_),
    .B1(_0419_),
    .B2(_2674_),
    .Y(_1422_));
 sky130_fd_sc_hd__a22o_1 _4641_ (.A1(\BitStream_buffer.BS_buffer[80] ),
    .A2(_2678_),
    .B1(_2681_),
    .B2(\BitStream_buffer.BS_buffer[81] ),
    .X(_1423_));
 sky130_fd_sc_hd__nor2_1 _4642_ (.A(_1422_),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__o22ai_1 _4643_ (.A1(_2757_),
    .A2(_2696_),
    .B1(_0440_),
    .B2(_2701_),
    .Y(_1425_));
 sky130_fd_sc_hd__a221oi_1 _4644_ (.A1(_2725_),
    .A2(_2688_),
    .B1(_2706_),
    .B2(_2692_),
    .C1(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__and4_1 _4645_ (.A(_1417_),
    .B(_1421_),
    .C(_1424_),
    .D(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__or2_1 _4646_ (.A(_2822_),
    .B(_2716_),
    .X(_1428_));
 sky130_fd_sc_hd__nand2_1 _4647_ (.A(_2719_),
    .B(_2820_),
    .Y(_1429_));
 sky130_fd_sc_hd__nand2_1 _4648_ (.A(_2723_),
    .B(_2804_),
    .Y(_1430_));
 sky130_fd_sc_hd__o2111a_1 _4649_ (.A1(_2795_),
    .A2(_2712_),
    .B1(_1428_),
    .C1(_1429_),
    .D1(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__o22ai_1 _4650_ (.A1(_2811_),
    .A2(_2734_),
    .B1(_0459_),
    .B2(_2738_),
    .Y(_1432_));
 sky130_fd_sc_hd__a221oi_1 _4651_ (.A1(_2792_),
    .A2(_2728_),
    .B1(\BitStream_buffer.BS_buffer[105] ),
    .B2(_2731_),
    .C1(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__nand2_1 _4652_ (.A(_2745_),
    .B(_2736_),
    .Y(_1434_));
 sky130_fd_sc_hd__nand2_1 _4653_ (.A(_2748_),
    .B(_2721_),
    .Y(_1435_));
 sky130_fd_sc_hd__or2_1 _4654_ (.A(_2733_),
    .B(_2752_),
    .X(_1436_));
 sky130_fd_sc_hd__o2111a_1 _4655_ (.A1(_2715_),
    .A2(_2743_),
    .B1(_1434_),
    .C1(_1435_),
    .D1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_2760_),
    .B(_2800_),
    .Y(_1438_));
 sky130_fd_sc_hd__nand2_1 _4657_ (.A(_2764_),
    .B(\BitStream_buffer.BS_buffer[94] ),
    .Y(_1439_));
 sky130_fd_sc_hd__or2_1 _4658_ (.A(_0568_),
    .B(_2770_),
    .X(_1440_));
 sky130_fd_sc_hd__o2111a_1 _4659_ (.A1(_2806_),
    .A2(_2758_),
    .B1(_1438_),
    .C1(_1439_),
    .D1(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__and4_1 _4660_ (.A(_1431_),
    .B(_1433_),
    .C(_1437_),
    .D(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__or2_1 _4661_ (.A(_2867_),
    .B(_2783_),
    .X(_1443_));
 sky130_fd_sc_hd__nand2_1 _4662_ (.A(_2786_),
    .B(\BitStream_buffer.BS_buffer[116] ),
    .Y(_1444_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_2790_),
    .B(\BitStream_buffer.BS_buffer[114] ),
    .Y(_1445_));
 sky130_fd_sc_hd__o2111a_1 _4664_ (.A1(_2894_),
    .A2(_2779_),
    .B1(_1443_),
    .C1(_1444_),
    .D1(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__nand2_1 _4665_ (.A(_2798_),
    .B(_2788_),
    .Y(_1447_));
 sky130_fd_sc_hd__nand2_1 _4666_ (.A(_2802_),
    .B(_2832_),
    .Y(_1448_));
 sky130_fd_sc_hd__or2_1 _4667_ (.A(_2782_),
    .B(_2807_),
    .X(_1449_));
 sky130_fd_sc_hd__o2111a_1 _4668_ (.A1(_2839_),
    .A2(_2796_),
    .B1(_1447_),
    .C1(_1448_),
    .D1(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__nand2_1 _4669_ (.A(_2814_),
    .B(\BitStream_buffer.BS_buffer[112] ),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_2818_),
    .B(_2836_),
    .Y(_1452_));
 sky130_fd_sc_hd__or2_1 _4671_ (.A(_2827_),
    .B(_2823_),
    .X(_1453_));
 sky130_fd_sc_hd__o2111a_1 _4672_ (.A1(_2898_),
    .A2(_2812_),
    .B1(_1451_),
    .C1(_1452_),
    .D1(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__nand2_1 _4673_ (.A(_2830_),
    .B(\BitStream_buffer.BS_buffer[118] ),
    .Y(_1455_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_2834_),
    .B(\BitStream_buffer.BS_buffer[120] ),
    .Y(_1456_));
 sky130_fd_sc_hd__or2_1 _4675_ (.A(_0601_),
    .B(_2840_),
    .X(_1457_));
 sky130_fd_sc_hd__o2111a_1 _4676_ (.A1(_2850_),
    .A2(_2828_),
    .B1(_1455_),
    .C1(_1456_),
    .D1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__and4_1 _4677_ (.A(_1446_),
    .B(_1450_),
    .C(_1454_),
    .D(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__or2_1 _4678_ (.A(_0638_),
    .B(_2851_),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _4679_ (.A(_2855_),
    .B(_0518_),
    .Y(_1461_));
 sky130_fd_sc_hd__nand2_1 _4680_ (.A(_2858_),
    .B(_3039_),
    .Y(_1462_));
 sky130_fd_sc_hd__o2111a_1 _4681_ (.A1(_0869_),
    .A2(_2848_),
    .B1(_1460_),
    .C1(_1461_),
    .D1(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__o22ai_1 _4682_ (.A1(_0604_),
    .A2(_2868_),
    .B1(_0476_),
    .B2(_2871_),
    .Y(_1464_));
 sky130_fd_sc_hd__a221oi_1 _4683_ (.A1(_0400_),
    .A2(_2862_),
    .B1(\BitStream_buffer.BS_buffer[1] ),
    .B2(_2866_),
    .C1(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__o22ai_1 _4684_ (.A1(_3024_),
    .A2(_2881_),
    .B1(_3027_),
    .B2(_2884_),
    .Y(_1466_));
 sky130_fd_sc_hd__a221oi_1 _4685_ (.A1(_0330_),
    .A2(_2875_),
    .B1(_0325_),
    .B2(_2879_),
    .C1(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(_2891_),
    .B(\BitStream_buffer.BS_buffer[124] ),
    .Y(_1468_));
 sky130_fd_sc_hd__or2_1 _4687_ (.A(_2880_),
    .B(_2895_),
    .X(_1469_));
 sky130_fd_sc_hd__or2_1 _4688_ (.A(_2845_),
    .B(_2899_),
    .X(_1470_));
 sky130_fd_sc_hd__o2111a_1 _4689_ (.A1(_0468_),
    .A2(_2889_),
    .B1(_1468_),
    .C1(_1469_),
    .D1(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__and4_1 _4690_ (.A(_1463_),
    .B(_1465_),
    .C(_1467_),
    .D(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__and4_1 _4691_ (.A(_1427_),
    .B(_1442_),
    .C(_1459_),
    .D(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__o22ai_1 _4692_ (.A1(_2939_),
    .A2(_2908_),
    .B1(_2942_),
    .B2(_2911_),
    .Y(_1474_));
 sky130_fd_sc_hd__o22ai_1 _4693_ (.A1(_0622_),
    .A2(_2915_),
    .B1(_0495_),
    .B2(_2919_),
    .Y(_1475_));
 sky130_fd_sc_hd__a22o_1 _4694_ (.A1(\BitStream_buffer.BS_buffer[48] ),
    .A2(_2923_),
    .B1(_2925_),
    .B2(\BitStream_buffer.BS_buffer[49] ),
    .X(_1476_));
 sky130_fd_sc_hd__a22o_1 _4695_ (.A1(\BitStream_buffer.BS_buffer[42] ),
    .A2(_2928_),
    .B1(_2930_),
    .B2(\BitStream_buffer.BS_buffer[43] ),
    .X(_1477_));
 sky130_fd_sc_hd__or4_1 _4696_ (.A(_1474_),
    .B(_1475_),
    .C(_1476_),
    .D(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__o22ai_1 _4697_ (.A1(_0858_),
    .A2(_2940_),
    .B1(_0750_),
    .B2(_2944_),
    .Y(_1479_));
 sky130_fd_sc_hd__a221oi_1 _4698_ (.A1(\BitStream_buffer.BS_buffer[54] ),
    .A2(_2934_),
    .B1(\BitStream_buffer.BS_buffer[55] ),
    .B2(_2937_),
    .C1(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__o22ai_1 _4699_ (.A1(_2963_),
    .A2(_2954_),
    .B1(_2968_),
    .B2(_2958_),
    .Y(_1481_));
 sky130_fd_sc_hd__a221oi_1 _4700_ (.A1(\BitStream_buffer.BS_buffer[50] ),
    .A2(_2948_),
    .B1(\BitStream_buffer.BS_buffer[51] ),
    .B2(_2951_),
    .C1(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__nand3b_1 _4701_ (.A_N(_1478_),
    .B(_1480_),
    .C(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__o22ai_1 _4702_ (.A1(_0508_),
    .A2(_2966_),
    .B1(_3009_),
    .B2(_2969_),
    .Y(_1484_));
 sky130_fd_sc_hd__o22ai_1 _4703_ (.A1(_0632_),
    .A2(_2973_),
    .B1(_0505_),
    .B2(_2976_),
    .Y(_1485_));
 sky130_fd_sc_hd__a22o_1 _4704_ (.A1(\BitStream_buffer.BS_buffer[64] ),
    .A2(_2980_),
    .B1(_2982_),
    .B2(\BitStream_buffer.BS_buffer[65] ),
    .X(_1486_));
 sky130_fd_sc_hd__a22o_1 _4705_ (.A1(\BitStream_buffer.BS_buffer[58] ),
    .A2(_2985_),
    .B1(_2987_),
    .B2(\BitStream_buffer.BS_buffer[59] ),
    .X(_1487_));
 sky130_fd_sc_hd__or4_1 _4706_ (.A(_1484_),
    .B(_1485_),
    .C(_1486_),
    .D(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__o22ai_1 _4707_ (.A1(_2664_),
    .A2(_2997_),
    .B1(_2671_),
    .B2(_3000_),
    .Y(_1489_));
 sky130_fd_sc_hd__a221oi_1 _4708_ (.A1(\BitStream_buffer.BS_buffer[66] ),
    .A2(_2991_),
    .B1(\BitStream_buffer.BS_buffer[67] ),
    .B2(_2994_),
    .C1(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__a2bb2o_1 _4709_ (.A1_N(_2631_),
    .A2_N(_3010_),
    .B1(\BitStream_buffer.BS_buffer[73] ),
    .B2(_3013_),
    .X(_1491_));
 sky130_fd_sc_hd__a221oi_1 _4710_ (.A1(\BitStream_buffer.BS_buffer[70] ),
    .A2(_3004_),
    .B1(\BitStream_buffer.BS_buffer[71] ),
    .B2(_3007_),
    .C1(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__nand3b_1 _4711_ (.A_N(_1488_),
    .B(_1490_),
    .C(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__nor2_1 _4712_ (.A(_3060_),
    .B(_3021_),
    .Y(_1494_));
 sky130_fd_sc_hd__o22ai_1 _4713_ (.A1(_0646_),
    .A2(_3025_),
    .B1(_0523_),
    .B2(_3029_),
    .Y(_1495_));
 sky130_fd_sc_hd__a22o_1 _4714_ (.A1(_0521_),
    .A2(_3033_),
    .B1(_3035_),
    .B2(\BitStream_buffer.BS_buffer[15] ),
    .X(_1496_));
 sky130_fd_sc_hd__a22o_1 _4715_ (.A1(_0770_),
    .A2(_3040_),
    .B1(_3042_),
    .B2(_3051_),
    .X(_1497_));
 sky130_fd_sc_hd__or4_1 _4716_ (.A(_1494_),
    .B(_1495_),
    .C(_1496_),
    .D(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__a22o_1 _4717_ (.A1(\BitStream_buffer.BS_buffer[22] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(\BitStream_buffer.BS_buffer[23] ),
    .X(_1499_));
 sky130_fd_sc_hd__o22ai_1 _4718_ (.A1(_0657_),
    .A2(_3054_),
    .B1(_0534_),
    .B2(_3057_),
    .Y(_1500_));
 sky130_fd_sc_hd__o22ai_1 _4719_ (.A1(_0660_),
    .A2(_3061_),
    .B1(_0537_),
    .B2(_0322_),
    .Y(_1501_));
 sky130_fd_sc_hd__a22o_1 _4720_ (.A1(\BitStream_buffer.BS_buffer[19] ),
    .A2(_0326_),
    .B1(_0328_),
    .B2(\BitStream_buffer.BS_buffer[18] ),
    .X(_1502_));
 sky130_fd_sc_hd__or4_1 _4721_ (.A(_1499_),
    .B(_1500_),
    .C(_1501_),
    .D(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__nor2_1 _4722_ (.A(_1498_),
    .B(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__o22ai_1 _4723_ (.A1(_2905_),
    .A2(_0343_),
    .B1(_2910_),
    .B2(_0346_),
    .Y(_1505_));
 sky130_fd_sc_hd__a221oi_1 _4724_ (.A1(\BitStream_buffer.BS_buffer[34] ),
    .A2(_0336_),
    .B1(\BitStream_buffer.BS_buffer[35] ),
    .B2(_0341_),
    .C1(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__o22ai_1 _4725_ (.A1(_0663_),
    .A2(_0356_),
    .B1(_0540_),
    .B2(_0359_),
    .Y(_1507_));
 sky130_fd_sc_hd__a221oi_1 _4726_ (.A1(_0387_),
    .A2(_0350_),
    .B1(\BitStream_buffer.BS_buffer[31] ),
    .B2(_0353_),
    .C1(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__o22ai_1 _4727_ (.A1(_0654_),
    .A2(_0371_),
    .B1(_0531_),
    .B2(_0374_),
    .Y(_1509_));
 sky130_fd_sc_hd__a221oi_1 _4728_ (.A1(\BitStream_buffer.BS_buffer[26] ),
    .A2(_0364_),
    .B1(\BitStream_buffer.BS_buffer[27] ),
    .B2(_0368_),
    .C1(_1509_),
    .Y(_1510_));
 sky130_fd_sc_hd__o22ai_1 _4729_ (.A1(_0847_),
    .A2(_0385_),
    .B1(_0739_),
    .B2(_0389_),
    .Y(_1511_));
 sky130_fd_sc_hd__a221oi_1 _4730_ (.A1(\BitStream_buffer.BS_buffer[38] ),
    .A2(_0378_),
    .B1(\BitStream_buffer.BS_buffer[39] ),
    .B2(_0383_),
    .C1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__and4_1 _4731_ (.A(_1506_),
    .B(_1508_),
    .C(_1510_),
    .D(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__nand2_1 _4732_ (.A(_1504_),
    .B(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__nor3_1 _4733_ (.A(_1483_),
    .B(_1493_),
    .C(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(_0398_),
    .B(_0527_),
    .Y(_1516_));
 sky130_fd_sc_hd__nand3_1 _4735_ (.A(_1473_),
    .B(_1515_),
    .C(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__inv_2 _4736_ (.A(\BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_1518_));
 sky130_fd_sc_hd__a21oi_1 _4737_ (.A1(_1518_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1519_));
 sky130_fd_sc_hd__o21a_1 _4738_ (.A1(_0672_),
    .A2(_1517_),
    .B1(_1519_),
    .X(_0311_));
 sky130_fd_sc_hd__o22ai_1 _4739_ (.A1(_0434_),
    .A2(_2629_),
    .B1(_2751_),
    .B2(_2636_),
    .Y(_1520_));
 sky130_fd_sc_hd__a221oi_1 _4740_ (.A1(_2768_),
    .A2(_2616_),
    .B1(_2762_),
    .B2(_2623_),
    .C1(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__nand2_1 _4741_ (.A(_2649_),
    .B(\BitStream_buffer.BS_buffer[77] ),
    .Y(_1522_));
 sky130_fd_sc_hd__or2_1 _4742_ (.A(_2698_),
    .B(_2655_),
    .X(_1523_));
 sky130_fd_sc_hd__or2_1 _4743_ (.A(_0419_),
    .B(_2660_),
    .X(_1524_));
 sky130_fd_sc_hd__o2111a_1 _4744_ (.A1(_0549_),
    .A2(_2645_),
    .B1(_1522_),
    .C1(_1523_),
    .D1(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__o22ai_1 _4745_ (.A1(_0686_),
    .A2(_2669_),
    .B1(_0560_),
    .B2(_2674_),
    .Y(_1526_));
 sky130_fd_sc_hd__a22o_1 _4746_ (.A1(\BitStream_buffer.BS_buffer[81] ),
    .A2(_2678_),
    .B1(_2681_),
    .B2(\BitStream_buffer.BS_buffer[82] ),
    .X(_1527_));
 sky130_fd_sc_hd__nor2_1 _4747_ (.A(_1526_),
    .B(_1527_),
    .Y(_1528_));
 sky130_fd_sc_hd__o22ai_1 _4748_ (.A1(_0437_),
    .A2(_2696_),
    .B1(_2757_),
    .B2(_2701_),
    .Y(_1529_));
 sky130_fd_sc_hd__a221oi_1 _4749_ (.A1(_2706_),
    .A2(_2688_),
    .B1(_2721_),
    .B2(_2692_),
    .C1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__and4_1 _4750_ (.A(_1521_),
    .B(_1525_),
    .C(_1528_),
    .D(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__or2_1 _4751_ (.A(_0459_),
    .B(_2716_),
    .X(_1532_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_2719_),
    .B(\BitStream_buffer.BS_buffer[101] ),
    .Y(_1533_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(_2723_),
    .B(\BitStream_buffer.BS_buffer[99] ),
    .Y(_1534_));
 sky130_fd_sc_hd__o2111a_1 _4754_ (.A1(_0450_),
    .A2(_2712_),
    .B1(_1532_),
    .C1(_1533_),
    .D1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__o22ai_1 _4755_ (.A1(_0456_),
    .A2(_2734_),
    .B1(_2811_),
    .B2(_2738_),
    .Y(_1536_));
 sky130_fd_sc_hd__a221oi_1 _4756_ (.A1(\BitStream_buffer.BS_buffer[105] ),
    .A2(_2728_),
    .B1(_2788_),
    .B2(_2731_),
    .C1(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_2745_),
    .B(\BitStream_buffer.BS_buffer[93] ),
    .Y(_1538_));
 sky130_fd_sc_hd__nand2_1 _4758_ (.A(_2748_),
    .B(_2714_),
    .Y(_1539_));
 sky130_fd_sc_hd__or2_1 _4759_ (.A(_0428_),
    .B(_2752_),
    .X(_1540_));
 sky130_fd_sc_hd__o2111a_1 _4760_ (.A1(_2737_),
    .A2(_2743_),
    .B1(_1538_),
    .C1(_1539_),
    .D1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__nand2_1 _4761_ (.A(_2760_),
    .B(\BitStream_buffer.BS_buffer[97] ),
    .Y(_1542_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(_2764_),
    .B(\BitStream_buffer.BS_buffer[95] ),
    .Y(_1543_));
 sky130_fd_sc_hd__or2_1 _4763_ (.A(_0694_),
    .B(_2770_),
    .X(_1544_));
 sky130_fd_sc_hd__o2111a_1 _4764_ (.A1(_0453_),
    .A2(_2758_),
    .B1(_1542_),
    .C1(_1543_),
    .D1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__and4_1 _4765_ (.A(_1535_),
    .B(_1537_),
    .C(_1541_),
    .D(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__or2_1 _4766_ (.A(_0473_),
    .B(_2783_),
    .X(_1547_));
 sky130_fd_sc_hd__nand2_1 _4767_ (.A(_2786_),
    .B(\BitStream_buffer.BS_buffer[117] ),
    .Y(_1548_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_2790_),
    .B(\BitStream_buffer.BS_buffer[115] ),
    .Y(_1549_));
 sky130_fd_sc_hd__o2111a_1 _4769_ (.A1(_2870_),
    .A2(_2779_),
    .B1(_1547_),
    .C1(_1548_),
    .D1(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__nand2_1 _4770_ (.A(_2798_),
    .B(_2781_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(_2802_),
    .B(_2838_),
    .Y(_1552_));
 sky130_fd_sc_hd__or2_1 _4772_ (.A(_0445_),
    .B(_2807_),
    .X(_1553_));
 sky130_fd_sc_hd__o2111a_1 _4773_ (.A1(_0464_),
    .A2(_2796_),
    .B1(_1551_),
    .C1(_1552_),
    .D1(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_2814_),
    .B(\BitStream_buffer.BS_buffer[113] ),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_1 _4775_ (.A(_2818_),
    .B(\BitStream_buffer.BS_buffer[111] ),
    .Y(_1556_));
 sky130_fd_sc_hd__or2_1 _4776_ (.A(_2888_),
    .B(_2823_),
    .X(_1557_));
 sky130_fd_sc_hd__o2111a_1 _4777_ (.A1(_0481_),
    .A2(_2812_),
    .B1(_1555_),
    .C1(_1556_),
    .D1(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__nand2_1 _4778_ (.A(_2830_),
    .B(\BitStream_buffer.BS_buffer[119] ),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(_2834_),
    .B(\BitStream_buffer.BS_buffer[121] ),
    .Y(_1560_));
 sky130_fd_sc_hd__or2_1 _4780_ (.A(_0727_),
    .B(_2840_),
    .X(_1561_));
 sky130_fd_sc_hd__o2111a_1 _4781_ (.A1(_0468_),
    .A2(_2828_),
    .B1(_1559_),
    .C1(_1560_),
    .D1(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__and4_1 _4782_ (.A(_1550_),
    .B(_1554_),
    .C(_1558_),
    .D(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__or2_1 _4783_ (.A(_0761_),
    .B(_2851_),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_1 _4784_ (.A(_2855_),
    .B(_3037_),
    .Y(_1565_));
 sky130_fd_sc_hd__nand2_1 _4785_ (.A(_2858_),
    .B(_3044_),
    .Y(_1566_));
 sky130_fd_sc_hd__o2111a_1 _4786_ (.A1(_3027_),
    .A2(_2848_),
    .B1(_1564_),
    .C1(_1565_),
    .D1(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__o22ai_1 _4787_ (.A1(_0730_),
    .A2(_2868_),
    .B1(_0604_),
    .B2(_2871_),
    .Y(_1568_));
 sky130_fd_sc_hd__a221oi_1 _4788_ (.A1(\BitStream_buffer.BS_buffer[1] ),
    .A2(_2862_),
    .B1(_3039_),
    .B2(_2865_),
    .C1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__o22ai_1 _4789_ (.A1(_0514_),
    .A2(_2881_),
    .B1(_3024_),
    .B2(_2884_),
    .Y(_1570_));
 sky130_fd_sc_hd__a221oi_1 _4790_ (.A1(_0325_),
    .A2(_2875_),
    .B1(_0527_),
    .B2(_2878_),
    .C1(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_1 _4791_ (.A(_2891_),
    .B(\BitStream_buffer.BS_buffer[125] ),
    .Y(_1572_));
 sky130_fd_sc_hd__or2_1 _4792_ (.A(_0476_),
    .B(_2895_),
    .X(_1573_));
 sky130_fd_sc_hd__or2_1 _4793_ (.A(_2883_),
    .B(_2899_),
    .X(_1574_));
 sky130_fd_sc_hd__o2111a_1 _4794_ (.A1(_2845_),
    .A2(_2889_),
    .B1(_1572_),
    .C1(_1573_),
    .D1(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__and4_1 _4795_ (.A(_1567_),
    .B(_1569_),
    .C(_1571_),
    .D(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__and4_1 _4796_ (.A(_1531_),
    .B(_1546_),
    .C(_1563_),
    .D(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__o22ai_1 _4797_ (.A1(_0492_),
    .A2(_2908_),
    .B1(_2939_),
    .B2(_2911_),
    .Y(_1578_));
 sky130_fd_sc_hd__o22ai_1 _4798_ (.A1(_2942_),
    .A2(_2915_),
    .B1(_0622_),
    .B2(_2919_),
    .Y(_1579_));
 sky130_fd_sc_hd__a22o_1 _4799_ (.A1(\BitStream_buffer.BS_buffer[49] ),
    .A2(_2923_),
    .B1(_2925_),
    .B2(\BitStream_buffer.BS_buffer[50] ),
    .X(_1580_));
 sky130_fd_sc_hd__a22o_1 _4800_ (.A1(\BitStream_buffer.BS_buffer[43] ),
    .A2(_2928_),
    .B1(_2930_),
    .B2(\BitStream_buffer.BS_buffer[44] ),
    .X(_1581_));
 sky130_fd_sc_hd__or4_1 _4801_ (.A(_1578_),
    .B(_1579_),
    .C(_1580_),
    .D(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__o22ai_1 _4802_ (.A1(_2999_),
    .A2(_2940_),
    .B1(_0858_),
    .B2(_2944_),
    .Y(_1583_));
 sky130_fd_sc_hd__a221oi_1 _4803_ (.A1(\BitStream_buffer.BS_buffer[55] ),
    .A2(_2934_),
    .B1(\BitStream_buffer.BS_buffer[56] ),
    .B2(_2937_),
    .C1(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__o22ai_1 _4804_ (.A1(_0499_),
    .A2(_2954_),
    .B1(_2963_),
    .B2(_2958_),
    .Y(_1585_));
 sky130_fd_sc_hd__a221oi_1 _4805_ (.A1(\BitStream_buffer.BS_buffer[51] ),
    .A2(_2948_),
    .B1(\BitStream_buffer.BS_buffer[52] ),
    .B2(_2951_),
    .C1(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__nand3b_1 _4806_ (.A_N(_1582_),
    .B(_1584_),
    .C(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__o22ai_1 _4807_ (.A1(_2640_),
    .A2(_2966_),
    .B1(_0508_),
    .B2(_2969_),
    .Y(_1588_));
 sky130_fd_sc_hd__o22ai_1 _4808_ (.A1(_3009_),
    .A2(_2973_),
    .B1(_0632_),
    .B2(_2976_),
    .Y(_1589_));
 sky130_fd_sc_hd__a22o_1 _4809_ (.A1(\BitStream_buffer.BS_buffer[65] ),
    .A2(_2980_),
    .B1(_2982_),
    .B2(\BitStream_buffer.BS_buffer[66] ),
    .X(_1590_));
 sky130_fd_sc_hd__a22o_1 _4810_ (.A1(\BitStream_buffer.BS_buffer[59] ),
    .A2(_2985_),
    .B1(_2987_),
    .B2(\BitStream_buffer.BS_buffer[60] ),
    .X(_1591_));
 sky130_fd_sc_hd__or4_1 _4811_ (.A(_1588_),
    .B(_1589_),
    .C(_1590_),
    .D(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__o22ai_1 _4812_ (.A1(_0415_),
    .A2(_2997_),
    .B1(_2664_),
    .B2(_3000_),
    .Y(_1593_));
 sky130_fd_sc_hd__a221oi_1 _4813_ (.A1(\BitStream_buffer.BS_buffer[67] ),
    .A2(_2991_),
    .B1(\BitStream_buffer.BS_buffer[68] ),
    .B2(_2994_),
    .C1(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__a2bb2o_1 _4814_ (.A1_N(_2625_),
    .A2_N(_3010_),
    .B1(\BitStream_buffer.BS_buffer[74] ),
    .B2(_3013_),
    .X(_1595_));
 sky130_fd_sc_hd__a221oi_1 _4815_ (.A1(\BitStream_buffer.BS_buffer[71] ),
    .A2(_3004_),
    .B1(\BitStream_buffer.BS_buffer[72] ),
    .B2(_3007_),
    .C1(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand3b_1 _4816_ (.A_N(_1592_),
    .B(_1594_),
    .C(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__nor2_1 _4817_ (.A(_0525_),
    .B(_3021_),
    .Y(_1598_));
 sky130_fd_sc_hd__o22ai_1 _4818_ (.A1(_0373_),
    .A2(_3025_),
    .B1(_0646_),
    .B2(_3029_),
    .Y(_1599_));
 sky130_fd_sc_hd__a22o_1 _4819_ (.A1(\BitStream_buffer.BS_buffer[15] ),
    .A2(_3033_),
    .B1(_3035_),
    .B2(_0363_),
    .X(_1600_));
 sky130_fd_sc_hd__a22o_1 _4820_ (.A1(_3051_),
    .A2(_3040_),
    .B1(_3042_),
    .B2(_0521_),
    .X(_1601_));
 sky130_fd_sc_hd__or4_1 _4821_ (.A(_1598_),
    .B(_1599_),
    .C(_1600_),
    .D(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__a22o_1 _4822_ (.A1(\BitStream_buffer.BS_buffer[23] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(\BitStream_buffer.BS_buffer[24] ),
    .X(_1603_));
 sky130_fd_sc_hd__o22ai_1 _4823_ (.A1(_0345_),
    .A2(_3054_),
    .B1(_0657_),
    .B2(_3057_),
    .Y(_1604_));
 sky130_fd_sc_hd__o22ai_1 _4824_ (.A1(_0358_),
    .A2(_3061_),
    .B1(_0660_),
    .B2(_0322_),
    .Y(_1605_));
 sky130_fd_sc_hd__a22o_1 _4825_ (.A1(\BitStream_buffer.BS_buffer[20] ),
    .A2(_0326_),
    .B1(_0328_),
    .B2(\BitStream_buffer.BS_buffer[19] ),
    .X(_1606_));
 sky130_fd_sc_hd__or4_1 _4826_ (.A(_1603_),
    .B(_1604_),
    .C(_1605_),
    .D(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__nor2_1 _4827_ (.A(_1602_),
    .B(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__o22ai_1 _4828_ (.A1(_0486_),
    .A2(_0343_),
    .B1(_2905_),
    .B2(_0346_),
    .Y(_1609_));
 sky130_fd_sc_hd__a221oi_1 _4829_ (.A1(\BitStream_buffer.BS_buffer[35] ),
    .A2(_0336_),
    .B1(\BitStream_buffer.BS_buffer[36] ),
    .B2(_0340_),
    .C1(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__o22ai_1 _4830_ (.A1(_2917_),
    .A2(_0356_),
    .B1(_0663_),
    .B2(_0359_),
    .Y(_1611_));
 sky130_fd_sc_hd__a221oi_1 _4831_ (.A1(\BitStream_buffer.BS_buffer[32] ),
    .A2(_0353_),
    .B1(\BitStream_buffer.BS_buffer[31] ),
    .B2(_0351_),
    .C1(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__o22ai_1 _4832_ (.A1(_0388_),
    .A2(_0371_),
    .B1(_0654_),
    .B2(_0374_),
    .Y(_1613_));
 sky130_fd_sc_hd__a221oi_1 _4833_ (.A1(\BitStream_buffer.BS_buffer[27] ),
    .A2(_0364_),
    .B1(\BitStream_buffer.BS_buffer[28] ),
    .B2(_0368_),
    .C1(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__o22ai_1 _4834_ (.A1(_2956_),
    .A2(_0385_),
    .B1(_0847_),
    .B2(_0389_),
    .Y(_1615_));
 sky130_fd_sc_hd__a221oi_1 _4835_ (.A1(\BitStream_buffer.BS_buffer[39] ),
    .A2(_0378_),
    .B1(\BitStream_buffer.BS_buffer[40] ),
    .B2(_0382_),
    .C1(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__and4_1 _4836_ (.A(_1610_),
    .B(_1612_),
    .C(_1614_),
    .D(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__nand2_1 _4837_ (.A(_1608_),
    .B(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__nor3_1 _4838_ (.A(_1587_),
    .B(_1597_),
    .C(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_0398_),
    .B(_0650_),
    .Y(_1620_));
 sky130_fd_sc_hd__nand3_1 _4840_ (.A(_1577_),
    .B(_1619_),
    .C(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__inv_2 _4841_ (.A(\BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_1622_));
 sky130_fd_sc_hd__a21oi_1 _4842_ (.A1(_1622_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1623_));
 sky130_fd_sc_hd__o21a_1 _4843_ (.A1(_0672_),
    .A2(_1621_),
    .B1(_1623_),
    .X(_0310_));
 sky130_fd_sc_hd__o22ai_1 _4844_ (.A1(_2769_),
    .A2(_2629_),
    .B1(_0434_),
    .B2(_2636_),
    .Y(_1624_));
 sky130_fd_sc_hd__a221oi_1 _4845_ (.A1(_2762_),
    .A2(_2616_),
    .B1(_2756_),
    .B2(_2623_),
    .C1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__nand2_1 _4846_ (.A(_2649_),
    .B(\BitStream_buffer.BS_buffer[78] ),
    .Y(_1626_));
 sky130_fd_sc_hd__or2_1 _4847_ (.A(_2694_),
    .B(_2655_),
    .X(_1627_));
 sky130_fd_sc_hd__or2_1 _4848_ (.A(_0560_),
    .B(_2660_),
    .X(_1628_));
 sky130_fd_sc_hd__o2111a_1 _4849_ (.A1(_2698_),
    .A2(_2645_),
    .B1(_1626_),
    .C1(_1627_),
    .D1(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__o22ai_1 _4850_ (.A1(_2742_),
    .A2(_2669_),
    .B1(_0686_),
    .B2(_2674_),
    .Y(_1630_));
 sky130_fd_sc_hd__a22o_1 _4851_ (.A1(\BitStream_buffer.BS_buffer[82] ),
    .A2(_2678_),
    .B1(_2681_),
    .B2(\BitStream_buffer.BS_buffer[83] ),
    .X(_1631_));
 sky130_fd_sc_hd__nor2_1 _4852_ (.A(_1630_),
    .B(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__o22ai_1 _4853_ (.A1(_2707_),
    .A2(_2696_),
    .B1(_0437_),
    .B2(_2701_),
    .Y(_1633_));
 sky130_fd_sc_hd__a221oi_1 _4854_ (.A1(_2721_),
    .A2(_2688_),
    .B1(_2714_),
    .B2(_2692_),
    .C1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__and4_1 _4855_ (.A(_1625_),
    .B(_1629_),
    .C(_1632_),
    .D(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__or2_1 _4856_ (.A(_2811_),
    .B(_2716_),
    .X(_1636_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(_2719_),
    .B(_2816_),
    .Y(_1637_));
 sky130_fd_sc_hd__nand2_1 _4858_ (.A(_2723_),
    .B(_2820_),
    .Y(_1638_));
 sky130_fd_sc_hd__o2111a_1 _4859_ (.A1(_2822_),
    .A2(_2712_),
    .B1(_1636_),
    .C1(_1637_),
    .D1(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__o22ai_1 _4860_ (.A1(_2775_),
    .A2(_2734_),
    .B1(_0456_),
    .B2(_2738_),
    .Y(_1640_));
 sky130_fd_sc_hd__a221oi_1 _4861_ (.A1(_2788_),
    .A2(_2728_),
    .B1(_2781_),
    .B2(_2731_),
    .C1(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _4862_ (.A(_2745_),
    .B(\BitStream_buffer.BS_buffer[94] ),
    .Y(_1642_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_2748_),
    .B(_2736_),
    .Y(_1643_));
 sky130_fd_sc_hd__or2_1 _4864_ (.A(_0568_),
    .B(_2752_),
    .X(_1644_));
 sky130_fd_sc_hd__o2111a_1 _4865_ (.A1(_2733_),
    .A2(_2743_),
    .B1(_1642_),
    .C1(_1643_),
    .D1(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__nand2_1 _4866_ (.A(_2760_),
    .B(_2804_),
    .Y(_1646_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(_2764_),
    .B(_2800_),
    .Y(_1647_));
 sky130_fd_sc_hd__or2_1 _4868_ (.A(_2806_),
    .B(_2770_),
    .X(_1648_));
 sky130_fd_sc_hd__o2111a_1 _4869_ (.A1(_2795_),
    .A2(_2758_),
    .B1(_1646_),
    .C1(_1647_),
    .D1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__and4_1 _4870_ (.A(_1639_),
    .B(_1641_),
    .C(_1645_),
    .D(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__or2_1 _4871_ (.A(_0601_),
    .B(_2783_),
    .X(_1651_));
 sky130_fd_sc_hd__nand2_1 _4872_ (.A(_2786_),
    .B(\BitStream_buffer.BS_buffer[118] ),
    .Y(_1652_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_2790_),
    .B(\BitStream_buffer.BS_buffer[116] ),
    .Y(_1653_));
 sky130_fd_sc_hd__o2111a_1 _4874_ (.A1(_2867_),
    .A2(_2779_),
    .B1(_1651_),
    .C1(_1652_),
    .D1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__nand2_1 _4875_ (.A(_2798_),
    .B(_2832_),
    .Y(_1655_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(_2802_),
    .B(_2836_),
    .Y(_1656_));
 sky130_fd_sc_hd__or2_1 _4877_ (.A(_2839_),
    .B(_2807_),
    .X(_1657_));
 sky130_fd_sc_hd__o2111a_1 _4878_ (.A1(_2827_),
    .A2(_2796_),
    .B1(_1655_),
    .C1(_1656_),
    .D1(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(_2814_),
    .B(\BitStream_buffer.BS_buffer[114] ),
    .Y(_1659_));
 sky130_fd_sc_hd__nand2_1 _4880_ (.A(_2818_),
    .B(\BitStream_buffer.BS_buffer[112] ),
    .Y(_1660_));
 sky130_fd_sc_hd__or2_1 _4881_ (.A(_2898_),
    .B(_2823_),
    .X(_1661_));
 sky130_fd_sc_hd__o2111a_1 _4882_ (.A1(_2894_),
    .A2(_2812_),
    .B1(_1659_),
    .C1(_1660_),
    .D1(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__nand2_1 _4883_ (.A(_2830_),
    .B(\BitStream_buffer.BS_buffer[120] ),
    .Y(_1663_));
 sky130_fd_sc_hd__nand2_1 _4884_ (.A(_2834_),
    .B(\BitStream_buffer.BS_buffer[122] ),
    .Y(_1664_));
 sky130_fd_sc_hd__or2_1 _4885_ (.A(_2850_),
    .B(_2840_),
    .X(_1665_));
 sky130_fd_sc_hd__o2111a_1 _4886_ (.A1(_2845_),
    .A2(_2828_),
    .B1(_1663_),
    .C1(_1664_),
    .D1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__and4_1 _4887_ (.A(_1654_),
    .B(_1658_),
    .C(_1662_),
    .D(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__or2_1 _4888_ (.A(_0869_),
    .B(_2851_),
    .X(_1668_));
 sky130_fd_sc_hd__nand2_1 _4889_ (.A(_2855_),
    .B(_0516_),
    .Y(_1669_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(_2858_),
    .B(_0518_),
    .Y(_1670_));
 sky130_fd_sc_hd__o2111a_1 _4891_ (.A1(_3024_),
    .A2(_2848_),
    .B1(_1668_),
    .C1(_1669_),
    .D1(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__o22ai_1 _4892_ (.A1(_3018_),
    .A2(_2868_),
    .B1(_0730_),
    .B2(_2871_),
    .Y(_1672_));
 sky130_fd_sc_hd__a221oi_1 _4893_ (.A1(_3039_),
    .A2(_2862_),
    .B1(_3044_),
    .B2(_2865_),
    .C1(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__o22ai_1 _4894_ (.A1(_0640_),
    .A2(_2881_),
    .B1(_0514_),
    .B2(_2884_),
    .Y(_1674_));
 sky130_fd_sc_hd__a221oi_1 _4895_ (.A1(_0527_),
    .A2(_2875_),
    .B1(_0650_),
    .B2(_2878_),
    .C1(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__nand2_1 _4896_ (.A(_2891_),
    .B(\BitStream_buffer.BS_buffer[126] ),
    .Y(_1676_));
 sky130_fd_sc_hd__or2_1 _4897_ (.A(_0604_),
    .B(_2895_),
    .X(_1677_));
 sky130_fd_sc_hd__or2_1 _4898_ (.A(_2880_),
    .B(_2899_),
    .X(_1678_));
 sky130_fd_sc_hd__o2111a_1 _4899_ (.A1(_2883_),
    .A2(_2889_),
    .B1(_1676_),
    .C1(_1677_),
    .D1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__and4_1 _4900_ (.A(_1671_),
    .B(_1673_),
    .C(_1675_),
    .D(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__and4_1 _4901_ (.A(_1635_),
    .B(_1650_),
    .C(_1667_),
    .D(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__o22ai_1 _4902_ (.A1(_0619_),
    .A2(_2908_),
    .B1(_0492_),
    .B2(_2911_),
    .Y(_1682_));
 sky130_fd_sc_hd__o22ai_1 _4903_ (.A1(_2939_),
    .A2(_2915_),
    .B1(_2942_),
    .B2(_2919_),
    .Y(_1683_));
 sky130_fd_sc_hd__a22o_1 _4904_ (.A1(\BitStream_buffer.BS_buffer[50] ),
    .A2(_2923_),
    .B1(_2925_),
    .B2(\BitStream_buffer.BS_buffer[51] ),
    .X(_1684_));
 sky130_fd_sc_hd__a22o_1 _4905_ (.A1(\BitStream_buffer.BS_buffer[44] ),
    .A2(_2928_),
    .B1(_2930_),
    .B2(\BitStream_buffer.BS_buffer[45] ),
    .X(_1685_));
 sky130_fd_sc_hd__or4_1 _4906_ (.A(_1682_),
    .B(_1683_),
    .C(_1684_),
    .D(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__o22ai_1 _4907_ (.A1(_2996_),
    .A2(_2940_),
    .B1(_2999_),
    .B2(_2944_),
    .Y(_1687_));
 sky130_fd_sc_hd__a221oi_1 _4908_ (.A1(\BitStream_buffer.BS_buffer[56] ),
    .A2(_2934_),
    .B1(\BitStream_buffer.BS_buffer[57] ),
    .B2(_2937_),
    .C1(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__o22ai_1 _4909_ (.A1(_0626_),
    .A2(_2954_),
    .B1(_0499_),
    .B2(_2958_),
    .Y(_1689_));
 sky130_fd_sc_hd__a221oi_1 _4910_ (.A1(\BitStream_buffer.BS_buffer[52] ),
    .A2(_2948_),
    .B1(\BitStream_buffer.BS_buffer[53] ),
    .B2(_2951_),
    .C1(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__nand3b_1 _4911_ (.A_N(_1686_),
    .B(_1688_),
    .C(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__o22ai_1 _4912_ (.A1(_2652_),
    .A2(_2966_),
    .B1(_2640_),
    .B2(_2969_),
    .Y(_1692_));
 sky130_fd_sc_hd__o22ai_1 _4913_ (.A1(_0508_),
    .A2(_2973_),
    .B1(_3009_),
    .B2(_2976_),
    .Y(_1693_));
 sky130_fd_sc_hd__a22o_1 _4914_ (.A1(\BitStream_buffer.BS_buffer[66] ),
    .A2(_2980_),
    .B1(_2982_),
    .B2(\BitStream_buffer.BS_buffer[67] ),
    .X(_1694_));
 sky130_fd_sc_hd__a22o_1 _4915_ (.A1(\BitStream_buffer.BS_buffer[60] ),
    .A2(_2985_),
    .B1(_2987_),
    .B2(\BitStream_buffer.BS_buffer[61] ),
    .X(_1695_));
 sky130_fd_sc_hd__or4_1 _4916_ (.A(_1692_),
    .B(_1693_),
    .C(_1694_),
    .D(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__o22ai_1 _4917_ (.A1(_0556_),
    .A2(_2997_),
    .B1(_0415_),
    .B2(_3000_),
    .Y(_1697_));
 sky130_fd_sc_hd__a221oi_1 _4918_ (.A1(\BitStream_buffer.BS_buffer[68] ),
    .A2(_2991_),
    .B1(\BitStream_buffer.BS_buffer[69] ),
    .B2(_2994_),
    .C1(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__a2bb2o_1 _4919_ (.A1_N(_0407_),
    .A2_N(_3010_),
    .B1(\BitStream_buffer.BS_buffer[75] ),
    .B2(_3013_),
    .X(_1699_));
 sky130_fd_sc_hd__a221oi_1 _4920_ (.A1(\BitStream_buffer.BS_buffer[72] ),
    .A2(_3004_),
    .B1(\BitStream_buffer.BS_buffer[73] ),
    .B2(_3007_),
    .C1(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand3b_1 _4921_ (.A_N(_1696_),
    .B(_1698_),
    .C(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__nor2_1 _4922_ (.A(_0648_),
    .B(_3021_),
    .Y(_1702_));
 sky130_fd_sc_hd__o22ai_1 _4923_ (.A1(_0370_),
    .A2(_3025_),
    .B1(_0373_),
    .B2(_3029_),
    .Y(_1703_));
 sky130_fd_sc_hd__a22o_1 _4924_ (.A1(_0363_),
    .A2(_3033_),
    .B1(_3035_),
    .B2(_0366_),
    .X(_1704_));
 sky130_fd_sc_hd__a22o_1 _4925_ (.A1(_0521_),
    .A2(_3040_),
    .B1(_3042_),
    .B2(\BitStream_buffer.BS_buffer[15] ),
    .X(_1705_));
 sky130_fd_sc_hd__or4_1 _4926_ (.A(_1702_),
    .B(_1703_),
    .C(_1704_),
    .D(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__a22o_1 _4927_ (.A1(\BitStream_buffer.BS_buffer[24] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(\BitStream_buffer.BS_buffer[25] ),
    .X(_1707_));
 sky130_fd_sc_hd__o22ai_1 _4928_ (.A1(_0342_),
    .A2(_3054_),
    .B1(_0345_),
    .B2(_3057_),
    .Y(_1708_));
 sky130_fd_sc_hd__o22ai_1 _4929_ (.A1(_0355_),
    .A2(_3061_),
    .B1(_0358_),
    .B2(_0322_),
    .Y(_1709_));
 sky130_fd_sc_hd__a22o_1 _4930_ (.A1(\BitStream_buffer.BS_buffer[21] ),
    .A2(_0326_),
    .B1(_0328_),
    .B2(\BitStream_buffer.BS_buffer[20] ),
    .X(_1710_));
 sky130_fd_sc_hd__or4_1 _4931_ (.A(_1707_),
    .B(_1708_),
    .C(_1709_),
    .D(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__nor2_1 _4932_ (.A(_1706_),
    .B(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__o22ai_1 _4933_ (.A1(_0613_),
    .A2(_0343_),
    .B1(_0486_),
    .B2(_0346_),
    .Y(_1713_));
 sky130_fd_sc_hd__a221oi_1 _4934_ (.A1(\BitStream_buffer.BS_buffer[36] ),
    .A2(_0336_),
    .B1(\BitStream_buffer.BS_buffer[37] ),
    .B2(_0340_),
    .C1(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__o22ai_1 _4935_ (.A1(_2914_),
    .A2(_0356_),
    .B1(_2917_),
    .B2(_0359_),
    .Y(_1715_));
 sky130_fd_sc_hd__a221oi_1 _4936_ (.A1(\BitStream_buffer.BS_buffer[32] ),
    .A2(_0350_),
    .B1(\BitStream_buffer.BS_buffer[33] ),
    .B2(_0353_),
    .C1(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__o22ai_1 _4937_ (.A1(_0384_),
    .A2(_0371_),
    .B1(_0388_),
    .B2(_0374_),
    .Y(_1717_));
 sky130_fd_sc_hd__a221oi_1 _4938_ (.A1(\BitStream_buffer.BS_buffer[28] ),
    .A2(_0364_),
    .B1(_0380_),
    .B2(_0368_),
    .C1(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__o22ai_1 _4939_ (.A1(_2953_),
    .A2(_0385_),
    .B1(_2956_),
    .B2(_0389_),
    .Y(_1719_));
 sky130_fd_sc_hd__a221oi_1 _4940_ (.A1(\BitStream_buffer.BS_buffer[40] ),
    .A2(_0378_),
    .B1(\BitStream_buffer.BS_buffer[41] ),
    .B2(_0382_),
    .C1(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__and4_1 _4941_ (.A(_1714_),
    .B(_1716_),
    .C(_1718_),
    .D(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(_1712_),
    .B(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__nor3_1 _4943_ (.A(_1691_),
    .B(_1701_),
    .C(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_1 _4944_ (.A(_0398_),
    .B(_0770_),
    .Y(_1724_));
 sky130_fd_sc_hd__nand3_1 _4945_ (.A(_1681_),
    .B(_1723_),
    .C(_1724_),
    .Y(_1725_));
 sky130_fd_sc_hd__inv_2 _4946_ (.A(\BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_1726_));
 sky130_fd_sc_hd__a21oi_1 _4947_ (.A1(_1726_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1727_));
 sky130_fd_sc_hd__o21a_1 _4948_ (.A1(_0672_),
    .A2(_1725_),
    .B1(_1727_),
    .X(_0309_));
 sky130_fd_sc_hd__o22ai_1 _4949_ (.A1(_0440_),
    .A2(_2629_),
    .B1(_2769_),
    .B2(_2636_),
    .Y(_1728_));
 sky130_fd_sc_hd__a221oi_1 _4950_ (.A1(_2756_),
    .A2(_2616_),
    .B1(_2725_),
    .B2(_2623_),
    .C1(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hd__nand2_1 _4951_ (.A(_2649_),
    .B(\BitStream_buffer.BS_buffer[79] ),
    .Y(_1730_));
 sky130_fd_sc_hd__or2_1 _4952_ (.A(_0419_),
    .B(_2655_),
    .X(_1731_));
 sky130_fd_sc_hd__or2_1 _4953_ (.A(_0686_),
    .B(_2660_),
    .X(_1732_));
 sky130_fd_sc_hd__o2111a_1 _4954_ (.A1(_2694_),
    .A2(_2645_),
    .B1(_1730_),
    .C1(_1731_),
    .D1(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__o22ai_1 _4955_ (.A1(_0431_),
    .A2(_2669_),
    .B1(_2742_),
    .B2(_2674_),
    .Y(_1734_));
 sky130_fd_sc_hd__a22o_1 _4956_ (.A1(\BitStream_buffer.BS_buffer[83] ),
    .A2(_2678_),
    .B1(_2681_),
    .B2(_2766_),
    .X(_1735_));
 sky130_fd_sc_hd__nor2_1 _4957_ (.A(_1734_),
    .B(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__o22ai_1 _4958_ (.A1(_0423_),
    .A2(_2696_),
    .B1(_2707_),
    .B2(_2701_),
    .Y(_1737_));
 sky130_fd_sc_hd__a221oi_1 _4959_ (.A1(_2714_),
    .A2(_2688_),
    .B1(_2736_),
    .B2(_2692_),
    .C1(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__and4_1 _4960_ (.A(_1729_),
    .B(_1733_),
    .C(_1736_),
    .D(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__or2_1 _4961_ (.A(_0456_),
    .B(_2716_),
    .X(_1740_));
 sky130_fd_sc_hd__nand2_1 _4962_ (.A(_2719_),
    .B(\BitStream_buffer.BS_buffer[103] ),
    .Y(_1741_));
 sky130_fd_sc_hd__nand2_1 _4963_ (.A(_2723_),
    .B(\BitStream_buffer.BS_buffer[101] ),
    .Y(_1742_));
 sky130_fd_sc_hd__o2111a_1 _4964_ (.A1(_0459_),
    .A2(_2712_),
    .B1(_1740_),
    .C1(_1741_),
    .D1(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__o22ai_1 _4965_ (.A1(_0444_),
    .A2(_2734_),
    .B1(_2775_),
    .B2(_2738_),
    .Y(_1744_));
 sky130_fd_sc_hd__a221oi_1 _4966_ (.A1(_2781_),
    .A2(_2728_),
    .B1(_2832_),
    .B2(_2731_),
    .C1(_1744_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2_1 _4967_ (.A(_2745_),
    .B(\BitStream_buffer.BS_buffer[95] ),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(_2748_),
    .B(\BitStream_buffer.BS_buffer[93] ),
    .Y(_1747_));
 sky130_fd_sc_hd__or2_1 _4969_ (.A(_0694_),
    .B(_2752_),
    .X(_1748_));
 sky130_fd_sc_hd__o2111a_1 _4970_ (.A1(_0428_),
    .A2(_2743_),
    .B1(_1746_),
    .C1(_1747_),
    .D1(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_2760_),
    .B(\BitStream_buffer.BS_buffer[99] ),
    .Y(_1750_));
 sky130_fd_sc_hd__nand2_1 _4972_ (.A(_2764_),
    .B(\BitStream_buffer.BS_buffer[97] ),
    .Y(_1751_));
 sky130_fd_sc_hd__or2_1 _4973_ (.A(_0453_),
    .B(_2770_),
    .X(_1752_));
 sky130_fd_sc_hd__o2111a_1 _4974_ (.A1(_0450_),
    .A2(_2758_),
    .B1(_1750_),
    .C1(_1751_),
    .D1(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__and4_1 _4975_ (.A(_1743_),
    .B(_1745_),
    .C(_1749_),
    .D(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__or2_1 _4976_ (.A(_0727_),
    .B(_2783_),
    .X(_1755_));
 sky130_fd_sc_hd__nand2_1 _4977_ (.A(_2786_),
    .B(\BitStream_buffer.BS_buffer[119] ),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(_2790_),
    .B(\BitStream_buffer.BS_buffer[117] ),
    .Y(_1757_));
 sky130_fd_sc_hd__o2111a_1 _4979_ (.A1(_0473_),
    .A2(_2779_),
    .B1(_1755_),
    .C1(_1756_),
    .D1(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__nand2_1 _4980_ (.A(_2798_),
    .B(_2838_),
    .Y(_1759_));
 sky130_fd_sc_hd__nand2_1 _4981_ (.A(_2802_),
    .B(\BitStream_buffer.BS_buffer[111] ),
    .Y(_1760_));
 sky130_fd_sc_hd__or2_1 _4982_ (.A(_0464_),
    .B(_2807_),
    .X(_1761_));
 sky130_fd_sc_hd__o2111a_1 _4983_ (.A1(_2888_),
    .A2(_2796_),
    .B1(_1759_),
    .C1(_1760_),
    .D1(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__nand2_1 _4984_ (.A(_2814_),
    .B(\BitStream_buffer.BS_buffer[115] ),
    .Y(_1763_));
 sky130_fd_sc_hd__nand2_1 _4985_ (.A(_2818_),
    .B(\BitStream_buffer.BS_buffer[113] ),
    .Y(_1764_));
 sky130_fd_sc_hd__or2_1 _4986_ (.A(_0481_),
    .B(_2823_),
    .X(_1765_));
 sky130_fd_sc_hd__o2111a_1 _4987_ (.A1(_2870_),
    .A2(_2812_),
    .B1(_1763_),
    .C1(_1764_),
    .D1(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_2830_),
    .B(\BitStream_buffer.BS_buffer[121] ),
    .Y(_1767_));
 sky130_fd_sc_hd__nand2_1 _4989_ (.A(_2834_),
    .B(\BitStream_buffer.BS_buffer[123] ),
    .Y(_1768_));
 sky130_fd_sc_hd__or2_1 _4990_ (.A(_0468_),
    .B(_2840_),
    .X(_1769_));
 sky130_fd_sc_hd__o2111a_1 _4991_ (.A1(_2883_),
    .A2(_2828_),
    .B1(_1767_),
    .C1(_1768_),
    .D1(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__and4_1 _4992_ (.A(_1758_),
    .B(_1762_),
    .C(_1766_),
    .D(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__or2_1 _4993_ (.A(_3027_),
    .B(_2851_),
    .X(_1772_));
 sky130_fd_sc_hd__nand2_1 _4994_ (.A(_2855_),
    .B(\BitStream_buffer.BS_buffer[7] ),
    .Y(_1773_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_2858_),
    .B(_3037_),
    .Y(_1774_));
 sky130_fd_sc_hd__o2111a_1 _4996_ (.A1(_0514_),
    .A2(_2848_),
    .B1(_1772_),
    .C1(_1773_),
    .D1(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__o22ai_1 _4997_ (.A1(_0512_),
    .A2(_2868_),
    .B1(_3018_),
    .B2(_2871_),
    .Y(_1776_));
 sky130_fd_sc_hd__a221oi_1 _4998_ (.A1(_3044_),
    .A2(_2862_),
    .B1(_0518_),
    .B2(_2865_),
    .C1(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__o22ai_1 _4999_ (.A1(_3063_),
    .A2(_2881_),
    .B1(_0640_),
    .B2(_2884_),
    .Y(_1778_));
 sky130_fd_sc_hd__a221oi_1 _5000_ (.A1(_0650_),
    .A2(_2875_),
    .B1(_0770_),
    .B2(_2878_),
    .C1(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__nand2_1 _5001_ (.A(_2891_),
    .B(\BitStream_buffer.BS_buffer[127] ),
    .Y(_1780_));
 sky130_fd_sc_hd__or2_1 _5002_ (.A(_0730_),
    .B(_2895_),
    .X(_1781_));
 sky130_fd_sc_hd__or2_1 _5003_ (.A(_0476_),
    .B(_2899_),
    .X(_1782_));
 sky130_fd_sc_hd__o2111a_1 _5004_ (.A1(_2880_),
    .A2(_2889_),
    .B1(_1780_),
    .C1(_1781_),
    .D1(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__and4_1 _5005_ (.A(_1775_),
    .B(_1777_),
    .C(_1779_),
    .D(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__and4_1 _5006_ (.A(_1739_),
    .B(_1754_),
    .C(_1771_),
    .D(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__o22ai_1 _5007_ (.A1(_2975_),
    .A2(_2908_),
    .B1(_0619_),
    .B2(_2911_),
    .Y(_1786_));
 sky130_fd_sc_hd__o22ai_1 _5008_ (.A1(_0492_),
    .A2(_2915_),
    .B1(_2939_),
    .B2(_2919_),
    .Y(_1787_));
 sky130_fd_sc_hd__a22o_1 _5009_ (.A1(\BitStream_buffer.BS_buffer[51] ),
    .A2(_2923_),
    .B1(_2925_),
    .B2(\BitStream_buffer.BS_buffer[52] ),
    .X(_1788_));
 sky130_fd_sc_hd__a22o_1 _5010_ (.A1(\BitStream_buffer.BS_buffer[45] ),
    .A2(_2928_),
    .B1(_2930_),
    .B2(\BitStream_buffer.BS_buffer[46] ),
    .X(_1789_));
 sky130_fd_sc_hd__or4_1 _5011_ (.A(_1786_),
    .B(_1787_),
    .C(_1788_),
    .D(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__o22ai_1 _5012_ (.A1(_0505_),
    .A2(_2940_),
    .B1(_2996_),
    .B2(_2944_),
    .Y(_1791_));
 sky130_fd_sc_hd__a221oi_1 _5013_ (.A1(\BitStream_buffer.BS_buffer[57] ),
    .A2(_2934_),
    .B1(\BitStream_buffer.BS_buffer[58] ),
    .B2(_2937_),
    .C1(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__o22ai_1 _5014_ (.A1(_0750_),
    .A2(_2954_),
    .B1(_0626_),
    .B2(_2958_),
    .Y(_1793_));
 sky130_fd_sc_hd__a221oi_1 _5015_ (.A1(\BitStream_buffer.BS_buffer[53] ),
    .A2(_2948_),
    .B1(\BitStream_buffer.BS_buffer[54] ),
    .B2(_2951_),
    .C1(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__nand3b_1 _5016_ (.A_N(_1790_),
    .B(_1792_),
    .C(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__o22ai_1 _5017_ (.A1(_0411_),
    .A2(_2966_),
    .B1(_2652_),
    .B2(_2969_),
    .Y(_1796_));
 sky130_fd_sc_hd__o22ai_1 _5018_ (.A1(_2640_),
    .A2(_2973_),
    .B1(_0508_),
    .B2(_2976_),
    .Y(_1797_));
 sky130_fd_sc_hd__a22o_1 _5019_ (.A1(\BitStream_buffer.BS_buffer[67] ),
    .A2(_2980_),
    .B1(_2982_),
    .B2(\BitStream_buffer.BS_buffer[68] ),
    .X(_1798_));
 sky130_fd_sc_hd__a22o_1 _5020_ (.A1(\BitStream_buffer.BS_buffer[61] ),
    .A2(_2985_),
    .B1(_2987_),
    .B2(\BitStream_buffer.BS_buffer[62] ),
    .X(_1799_));
 sky130_fd_sc_hd__or4_1 _5021_ (.A(_1796_),
    .B(_1797_),
    .C(_1798_),
    .D(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__o22ai_1 _5022_ (.A1(_2631_),
    .A2(_2997_),
    .B1(_0556_),
    .B2(_3000_),
    .Y(_1801_));
 sky130_fd_sc_hd__a221oi_1 _5023_ (.A1(\BitStream_buffer.BS_buffer[69] ),
    .A2(_2991_),
    .B1(\BitStream_buffer.BS_buffer[70] ),
    .B2(_2994_),
    .C1(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__a2bb2o_1 _5024_ (.A1_N(_0549_),
    .A2_N(_3010_),
    .B1(\BitStream_buffer.BS_buffer[76] ),
    .B2(_3013_),
    .X(_1803_));
 sky130_fd_sc_hd__a221oi_1 _5025_ (.A1(\BitStream_buffer.BS_buffer[73] ),
    .A2(_3004_),
    .B1(\BitStream_buffer.BS_buffer[74] ),
    .B2(_3007_),
    .C1(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__nand3b_1 _5026_ (.A_N(_1800_),
    .B(_1802_),
    .C(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__nor2_1 _5027_ (.A(_3056_),
    .B(_3021_),
    .Y(_1806_));
 sky130_fd_sc_hd__o22ai_1 _5028_ (.A1(_0537_),
    .A2(_3025_),
    .B1(_0370_),
    .B2(_3029_),
    .Y(_1807_));
 sky130_fd_sc_hd__a22o_1 _5029_ (.A1(_0366_),
    .A2(_3033_),
    .B1(_3035_),
    .B2(\BitStream_buffer.BS_buffer[18] ),
    .X(_1808_));
 sky130_fd_sc_hd__a22o_1 _5030_ (.A1(\BitStream_buffer.BS_buffer[15] ),
    .A2(_3040_),
    .B1(_3042_),
    .B2(_0363_),
    .X(_1809_));
 sky130_fd_sc_hd__or4_1 _5031_ (.A(_1806_),
    .B(_1807_),
    .C(_1808_),
    .D(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__a22o_1 _5032_ (.A1(\BitStream_buffer.BS_buffer[25] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(\BitStream_buffer.BS_buffer[26] ),
    .X(_1811_));
 sky130_fd_sc_hd__o22ai_1 _5033_ (.A1(_0531_),
    .A2(_3054_),
    .B1(_0342_),
    .B2(_3057_),
    .Y(_1812_));
 sky130_fd_sc_hd__o22ai_1 _5034_ (.A1(_0534_),
    .A2(_3061_),
    .B1(_0355_),
    .B2(_0322_),
    .Y(_1813_));
 sky130_fd_sc_hd__a22o_1 _5035_ (.A1(\BitStream_buffer.BS_buffer[22] ),
    .A2(_0326_),
    .B1(_0328_),
    .B2(\BitStream_buffer.BS_buffer[21] ),
    .X(_1814_));
 sky130_fd_sc_hd__or4_1 _5036_ (.A(_1811_),
    .B(_1812_),
    .C(_1813_),
    .D(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__nor2_1 _5037_ (.A(_1810_),
    .B(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__o22ai_1 _5038_ (.A1(_0739_),
    .A2(_0343_),
    .B1(_0613_),
    .B2(_0346_),
    .Y(_1817_));
 sky130_fd_sc_hd__a221oi_1 _5039_ (.A1(\BitStream_buffer.BS_buffer[37] ),
    .A2(_0336_),
    .B1(\BitStream_buffer.BS_buffer[38] ),
    .B2(_0340_),
    .C1(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__o22ai_1 _5040_ (.A1(_2910_),
    .A2(_0356_),
    .B1(_2914_),
    .B2(_0359_),
    .Y(_1819_));
 sky130_fd_sc_hd__a221oi_1 _5041_ (.A1(\BitStream_buffer.BS_buffer[33] ),
    .A2(_0350_),
    .B1(\BitStream_buffer.BS_buffer[34] ),
    .B2(_0353_),
    .C1(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__o22ai_1 _5042_ (.A1(_0540_),
    .A2(_0371_),
    .B1(_0384_),
    .B2(_0374_),
    .Y(_1821_));
 sky130_fd_sc_hd__a221oi_1 _5043_ (.A1(_0380_),
    .A2(_0364_),
    .B1(_0387_),
    .B2(_0368_),
    .C1(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__o22ai_1 _5044_ (.A1(_0495_),
    .A2(_0385_),
    .B1(_2953_),
    .B2(_0389_),
    .Y(_1823_));
 sky130_fd_sc_hd__a221oi_1 _5045_ (.A1(\BitStream_buffer.BS_buffer[41] ),
    .A2(_0378_),
    .B1(\BitStream_buffer.BS_buffer[42] ),
    .B2(_0382_),
    .C1(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__and4_1 _5046_ (.A(_1818_),
    .B(_1820_),
    .C(_1822_),
    .D(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__nand2_1 _5047_ (.A(_1816_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__nor3_1 _5048_ (.A(_1795_),
    .B(_1805_),
    .C(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_0398_),
    .B(_3051_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand3_1 _5050_ (.A(_1785_),
    .B(_1827_),
    .C(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__inv_2 _5051_ (.A(\BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_1830_));
 sky130_fd_sc_hd__a21oi_1 _5052_ (.A1(_1830_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1831_));
 sky130_fd_sc_hd__o21a_1 _5053_ (.A1(_0672_),
    .A2(_1829_),
    .B1(_1831_),
    .X(_0308_));
 sky130_fd_sc_hd__o22ai_1 _5054_ (.A1(_2757_),
    .A2(_2629_),
    .B1(_0440_),
    .B2(_2636_),
    .Y(_1832_));
 sky130_fd_sc_hd__a221oi_1 _5055_ (.A1(_2725_),
    .A2(_2616_),
    .B1(_2706_),
    .B2(_2623_),
    .C1(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _5056_ (.A(_2649_),
    .B(\BitStream_buffer.BS_buffer[80] ),
    .Y(_1834_));
 sky130_fd_sc_hd__or2_1 _5057_ (.A(_0560_),
    .B(_2655_),
    .X(_1835_));
 sky130_fd_sc_hd__or2_1 _5058_ (.A(_2742_),
    .B(_2660_),
    .X(_1836_));
 sky130_fd_sc_hd__o2111a_1 _5059_ (.A1(_0419_),
    .A2(_2645_),
    .B1(_1834_),
    .C1(_1835_),
    .D1(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__o22ai_1 _5060_ (.A1(_2751_),
    .A2(_2669_),
    .B1(_0431_),
    .B2(_2674_),
    .Y(_1838_));
 sky130_fd_sc_hd__a22o_1 _5061_ (.A1(_2766_),
    .A2(_2678_),
    .B1(_2681_),
    .B2(_2768_),
    .X(_1839_));
 sky130_fd_sc_hd__nor2_1 _5062_ (.A(_1838_),
    .B(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__o22ai_1 _5063_ (.A1(_2715_),
    .A2(_2696_),
    .B1(_0423_),
    .B2(_2701_),
    .Y(_1841_));
 sky130_fd_sc_hd__a221oi_1 _5064_ (.A1(_2736_),
    .A2(_2688_),
    .B1(\BitStream_buffer.BS_buffer[93] ),
    .B2(_2692_),
    .C1(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__and4_1 _5065_ (.A(_1833_),
    .B(_1837_),
    .C(_1840_),
    .D(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__or2_1 _5066_ (.A(_2775_),
    .B(_2716_),
    .X(_1844_));
 sky130_fd_sc_hd__nand2_1 _5067_ (.A(_2719_),
    .B(_2792_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2_1 _5068_ (.A(_2723_),
    .B(_2816_),
    .Y(_1846_));
 sky130_fd_sc_hd__o2111a_1 _5069_ (.A1(_2811_),
    .A2(_2712_),
    .B1(_1844_),
    .C1(_1845_),
    .D1(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__o22ai_1 _5070_ (.A1(_2782_),
    .A2(_2734_),
    .B1(_0444_),
    .B2(_2738_),
    .Y(_1848_));
 sky130_fd_sc_hd__a221oi_1 _5071_ (.A1(_2832_),
    .A2(_2728_),
    .B1(_2838_),
    .B2(_2731_),
    .C1(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__nand2_1 _5072_ (.A(_2745_),
    .B(_2800_),
    .Y(_1850_));
 sky130_fd_sc_hd__nand2_1 _5073_ (.A(_2748_),
    .B(\BitStream_buffer.BS_buffer[94] ),
    .Y(_1851_));
 sky130_fd_sc_hd__or2_1 _5074_ (.A(_2806_),
    .B(_2752_),
    .X(_1852_));
 sky130_fd_sc_hd__o2111a_1 _5075_ (.A1(_0568_),
    .A2(_2743_),
    .B1(_1850_),
    .C1(_1851_),
    .D1(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__nand2_1 _5076_ (.A(_2760_),
    .B(_2820_),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _5077_ (.A(_2764_),
    .B(_2804_),
    .Y(_1855_));
 sky130_fd_sc_hd__or2_1 _5078_ (.A(_2795_),
    .B(_2770_),
    .X(_1856_));
 sky130_fd_sc_hd__o2111a_1 _5079_ (.A1(_2822_),
    .A2(_2758_),
    .B1(_1854_),
    .C1(_1855_),
    .D1(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__and4_1 _5080_ (.A(_1847_),
    .B(_1849_),
    .C(_1853_),
    .D(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__or2_1 _5081_ (.A(_2850_),
    .B(_2783_),
    .X(_1859_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_2786_),
    .B(\BitStream_buffer.BS_buffer[120] ),
    .Y(_1860_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_2790_),
    .B(\BitStream_buffer.BS_buffer[118] ),
    .Y(_1861_));
 sky130_fd_sc_hd__o2111a_1 _5084_ (.A1(_0601_),
    .A2(_2779_),
    .B1(_1859_),
    .C1(_1860_),
    .D1(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_2798_),
    .B(_2836_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_2802_),
    .B(\BitStream_buffer.BS_buffer[112] ),
    .Y(_1864_));
 sky130_fd_sc_hd__or2_1 _5087_ (.A(_2827_),
    .B(_2807_),
    .X(_1865_));
 sky130_fd_sc_hd__o2111a_1 _5088_ (.A1(_2898_),
    .A2(_2796_),
    .B1(_1863_),
    .C1(_1864_),
    .D1(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__nand2_1 _5089_ (.A(_2814_),
    .B(\BitStream_buffer.BS_buffer[116] ),
    .Y(_1867_));
 sky130_fd_sc_hd__nand2_1 _5090_ (.A(_2818_),
    .B(\BitStream_buffer.BS_buffer[114] ),
    .Y(_1868_));
 sky130_fd_sc_hd__or2_1 _5091_ (.A(_2894_),
    .B(_2823_),
    .X(_1869_));
 sky130_fd_sc_hd__o2111a_1 _5092_ (.A1(_2867_),
    .A2(_2812_),
    .B1(_1867_),
    .C1(_1868_),
    .D1(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__nand2_1 _5093_ (.A(_2830_),
    .B(\BitStream_buffer.BS_buffer[122] ),
    .Y(_1871_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_2834_),
    .B(\BitStream_buffer.BS_buffer[124] ),
    .Y(_1872_));
 sky130_fd_sc_hd__or2_1 _5095_ (.A(_2845_),
    .B(_2840_),
    .X(_1873_));
 sky130_fd_sc_hd__o2111a_1 _5096_ (.A1(_2880_),
    .A2(_2828_),
    .B1(_1871_),
    .C1(_1872_),
    .D1(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__and4_1 _5097_ (.A(_1862_),
    .B(_1866_),
    .C(_1870_),
    .D(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__or2_1 _5098_ (.A(_3024_),
    .B(_2851_),
    .X(_1876_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_2855_),
    .B(_0330_),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _5100_ (.A(_2858_),
    .B(_0516_),
    .Y(_1878_));
 sky130_fd_sc_hd__o2111a_1 _5101_ (.A1(_0640_),
    .A2(_2848_),
    .B1(_1876_),
    .C1(_1877_),
    .D1(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__o22ai_1 _5102_ (.A1(_0638_),
    .A2(_2868_),
    .B1(_0512_),
    .B2(_2871_),
    .Y(_1880_));
 sky130_fd_sc_hd__a221oi_1 _5103_ (.A1(_0518_),
    .A2(_2862_),
    .B1(_3037_),
    .B2(_2865_),
    .C1(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hd__o22ai_1 _5104_ (.A1(_3060_),
    .A2(_2881_),
    .B1(_3063_),
    .B2(_2884_),
    .Y(_1882_));
 sky130_fd_sc_hd__a221oi_1 _5105_ (.A1(_0770_),
    .A2(_2875_),
    .B1(_3051_),
    .B2(_2878_),
    .C1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__nand2_1 _5106_ (.A(_2891_),
    .B(_0400_),
    .Y(_1884_));
 sky130_fd_sc_hd__or2_1 _5107_ (.A(_3018_),
    .B(_2895_),
    .X(_1885_));
 sky130_fd_sc_hd__or2_1 _5108_ (.A(_0604_),
    .B(_2899_),
    .X(_1886_));
 sky130_fd_sc_hd__o2111a_1 _5109_ (.A1(_0476_),
    .A2(_2889_),
    .B1(_1884_),
    .C1(_1885_),
    .D1(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__and4_1 _5110_ (.A(_1879_),
    .B(_1881_),
    .C(_1883_),
    .D(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__and4_1 _5111_ (.A(_1843_),
    .B(_1858_),
    .C(_1875_),
    .D(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__o22ai_1 _5112_ (.A1(_2972_),
    .A2(_2908_),
    .B1(_2975_),
    .B2(_2911_),
    .Y(_1890_));
 sky130_fd_sc_hd__o22ai_1 _5113_ (.A1(_0619_),
    .A2(_2915_),
    .B1(_0492_),
    .B2(_2919_),
    .Y(_1891_));
 sky130_fd_sc_hd__a22o_1 _5114_ (.A1(\BitStream_buffer.BS_buffer[52] ),
    .A2(_2923_),
    .B1(_2925_),
    .B2(\BitStream_buffer.BS_buffer[53] ),
    .X(_1892_));
 sky130_fd_sc_hd__a22o_1 _5115_ (.A1(\BitStream_buffer.BS_buffer[46] ),
    .A2(_2928_),
    .B1(_2930_),
    .B2(\BitStream_buffer.BS_buffer[47] ),
    .X(_1893_));
 sky130_fd_sc_hd__or4_1 _5116_ (.A(_1890_),
    .B(_1891_),
    .C(_1892_),
    .D(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__o22ai_1 _5117_ (.A1(_0632_),
    .A2(_2940_),
    .B1(_0505_),
    .B2(_2944_),
    .Y(_1895_));
 sky130_fd_sc_hd__a221oi_1 _5118_ (.A1(\BitStream_buffer.BS_buffer[58] ),
    .A2(_2934_),
    .B1(\BitStream_buffer.BS_buffer[59] ),
    .B2(_2937_),
    .C1(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__o22ai_1 _5119_ (.A1(_0858_),
    .A2(_2954_),
    .B1(_0750_),
    .B2(_2958_),
    .Y(_1897_));
 sky130_fd_sc_hd__a221oi_1 _5120_ (.A1(\BitStream_buffer.BS_buffer[54] ),
    .A2(_2948_),
    .B1(\BitStream_buffer.BS_buffer[55] ),
    .B2(_2951_),
    .C1(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__nand3b_1 _5121_ (.A_N(_1894_),
    .B(_1896_),
    .C(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__o22ai_1 _5122_ (.A1(_2658_),
    .A2(_2966_),
    .B1(_0411_),
    .B2(_2969_),
    .Y(_1900_));
 sky130_fd_sc_hd__o22ai_1 _5123_ (.A1(_2652_),
    .A2(_2973_),
    .B1(_2640_),
    .B2(_2976_),
    .Y(_1901_));
 sky130_fd_sc_hd__a22o_1 _5124_ (.A1(\BitStream_buffer.BS_buffer[68] ),
    .A2(_2980_),
    .B1(_2982_),
    .B2(\BitStream_buffer.BS_buffer[69] ),
    .X(_1902_));
 sky130_fd_sc_hd__a22o_1 _5125_ (.A1(\BitStream_buffer.BS_buffer[62] ),
    .A2(_2985_),
    .B1(_2987_),
    .B2(\BitStream_buffer.BS_buffer[63] ),
    .X(_1903_));
 sky130_fd_sc_hd__or4_1 _5126_ (.A(_1900_),
    .B(_1901_),
    .C(_1902_),
    .D(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__o22ai_1 _5127_ (.A1(_2625_),
    .A2(_2997_),
    .B1(_2631_),
    .B2(_3000_),
    .Y(_1905_));
 sky130_fd_sc_hd__a221oi_1 _5128_ (.A1(\BitStream_buffer.BS_buffer[70] ),
    .A2(_2991_),
    .B1(\BitStream_buffer.BS_buffer[71] ),
    .B2(_2994_),
    .C1(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__a2bb2o_1 _5129_ (.A1_N(_2698_),
    .A2_N(_3010_),
    .B1(\BitStream_buffer.BS_buffer[77] ),
    .B2(_3013_),
    .X(_1907_));
 sky130_fd_sc_hd__a221oi_1 _5130_ (.A1(\BitStream_buffer.BS_buffer[74] ),
    .A2(_3004_),
    .B1(\BitStream_buffer.BS_buffer[75] ),
    .B2(_3007_),
    .C1(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__nand3b_1 _5131_ (.A_N(_1904_),
    .B(_1906_),
    .C(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__nor2_1 _5132_ (.A(_3053_),
    .B(_3021_),
    .Y(_1910_));
 sky130_fd_sc_hd__o22ai_1 _5133_ (.A1(_0660_),
    .A2(_3025_),
    .B1(_0537_),
    .B2(_3029_),
    .Y(_1911_));
 sky130_fd_sc_hd__a22o_1 _5134_ (.A1(\BitStream_buffer.BS_buffer[18] ),
    .A2(_3033_),
    .B1(_3035_),
    .B2(\BitStream_buffer.BS_buffer[19] ),
    .X(_1912_));
 sky130_fd_sc_hd__a22o_1 _5135_ (.A1(_0363_),
    .A2(_3040_),
    .B1(_3042_),
    .B2(_0366_),
    .X(_1913_));
 sky130_fd_sc_hd__or4_1 _5136_ (.A(_1910_),
    .B(_1911_),
    .C(_1912_),
    .D(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__a22o_1 _5137_ (.A1(\BitStream_buffer.BS_buffer[26] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(\BitStream_buffer.BS_buffer[27] ),
    .X(_1915_));
 sky130_fd_sc_hd__o22ai_1 _5138_ (.A1(_0654_),
    .A2(_3054_),
    .B1(_0531_),
    .B2(_3057_),
    .Y(_1916_));
 sky130_fd_sc_hd__o22ai_1 _5139_ (.A1(_0657_),
    .A2(_3061_),
    .B1(_0534_),
    .B2(_0322_),
    .Y(_1917_));
 sky130_fd_sc_hd__a22o_1 _5140_ (.A1(\BitStream_buffer.BS_buffer[23] ),
    .A2(_0326_),
    .B1(_0328_),
    .B2(\BitStream_buffer.BS_buffer[22] ),
    .X(_1918_));
 sky130_fd_sc_hd__or4_1 _5141_ (.A(_1915_),
    .B(_1916_),
    .C(_1917_),
    .D(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__nor2_1 _5142_ (.A(_1914_),
    .B(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__o22ai_1 _5143_ (.A1(_0847_),
    .A2(_0343_),
    .B1(_0739_),
    .B2(_0346_),
    .Y(_1921_));
 sky130_fd_sc_hd__a221oi_1 _5144_ (.A1(\BitStream_buffer.BS_buffer[38] ),
    .A2(_0336_),
    .B1(\BitStream_buffer.BS_buffer[39] ),
    .B2(_0340_),
    .C1(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__o22ai_1 _5145_ (.A1(_2905_),
    .A2(_0356_),
    .B1(_2910_),
    .B2(_0359_),
    .Y(_1923_));
 sky130_fd_sc_hd__a221oi_1 _5146_ (.A1(\BitStream_buffer.BS_buffer[34] ),
    .A2(_0350_),
    .B1(\BitStream_buffer.BS_buffer[35] ),
    .B2(_0353_),
    .C1(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__o22ai_1 _5147_ (.A1(_0663_),
    .A2(_0371_),
    .B1(_0540_),
    .B2(_0374_),
    .Y(_1925_));
 sky130_fd_sc_hd__a221oi_1 _5148_ (.A1(_0387_),
    .A2(_0364_),
    .B1(\BitStream_buffer.BS_buffer[31] ),
    .B2(_0368_),
    .C1(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__o22ai_1 _5149_ (.A1(_0622_),
    .A2(_0385_),
    .B1(_0495_),
    .B2(_0389_),
    .Y(_1927_));
 sky130_fd_sc_hd__a221oi_1 _5150_ (.A1(\BitStream_buffer.BS_buffer[42] ),
    .A2(_0378_),
    .B1(\BitStream_buffer.BS_buffer[43] ),
    .B2(_0382_),
    .C1(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__and4_1 _5151_ (.A(_1922_),
    .B(_1924_),
    .C(_1926_),
    .D(_1928_),
    .X(_1929_));
 sky130_fd_sc_hd__nand2_1 _5152_ (.A(_1920_),
    .B(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__nor3_1 _5153_ (.A(_1899_),
    .B(_1909_),
    .C(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _5154_ (.A(_0398_),
    .B(_0521_),
    .Y(_1932_));
 sky130_fd_sc_hd__nand3_1 _5155_ (.A(_1889_),
    .B(_1931_),
    .C(_1932_),
    .Y(_1933_));
 sky130_fd_sc_hd__inv_2 _5156_ (.A(\BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_1934_));
 sky130_fd_sc_hd__a21oi_1 _5157_ (.A1(_1934_),
    .A2(_2598_),
    .B1(_0674_),
    .Y(_1935_));
 sky130_fd_sc_hd__o21a_1 _5158_ (.A1(_0672_),
    .A2(_1933_),
    .B1(_1935_),
    .X(_0307_));
 sky130_fd_sc_hd__inv_2 _5159_ (.A(net34),
    .Y(_1936_));
 sky130_fd_sc_hd__nor2_1 _5160_ (.A(net33),
    .B(net32),
    .Y(_1937_));
 sky130_fd_sc_hd__nor2_2 _5161_ (.A(_1936_),
    .B(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__and2_1 _5162_ (.A(_1937_),
    .B(_1936_),
    .X(_1939_));
 sky130_fd_sc_hd__nor2_1 _5163_ (.A(net30),
    .B(net29),
    .Y(_1940_));
 sky130_fd_sc_hd__inv_2 _5164_ (.A(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__nand2_1 _5165_ (.A(net198),
    .B(net29),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5166_ (.A(_1941_),
    .B(net199),
    .Y(_1943_));
 sky130_fd_sc_hd__o21ai_4 _5167_ (.A1(_1938_),
    .A2(_1939_),
    .B1(net200),
    .Y(_1944_));
 sky130_fd_sc_hd__inv_2 _5168_ (.A(\BitStream_buffer.buffer_index[6] ),
    .Y(_1945_));
 sky130_fd_sc_hd__inv_2 _5169_ (.A(\BitStream_buffer.buffer_index[5] ),
    .Y(_1946_));
 sky130_fd_sc_hd__inv_2 _5170_ (.A(\BitStream_buffer.buffer_index[4] ),
    .Y(_1947_));
 sky130_fd_sc_hd__and3_1 _5171_ (.A(_1945_),
    .B(_1946_),
    .C(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__nand2_4 _5172_ (.A(_1944_),
    .B(_1948_),
    .Y(_1949_));
 sky130_fd_sc_hd__clkbuf_4 _5173_ (.A(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__mux2_1 _5174_ (.A0(net7),
    .A1(_0400_),
    .S(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__clkbuf_2 _5175_ (.A(_0404_),
    .X(_1952_));
 sky130_fd_sc_hd__and2_1 _5176_ (.A(_1951_),
    .B(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__clkbuf_1 _5177_ (.A(_1953_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _5178_ (.A0(net6),
    .A1(\BitStream_buffer.BS_buffer[1] ),
    .S(_1950_),
    .X(_1954_));
 sky130_fd_sc_hd__and2_1 _5179_ (.A(_1954_),
    .B(_1952_),
    .X(_1955_));
 sky130_fd_sc_hd__clkbuf_1 _5180_ (.A(_1955_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _5181_ (.A0(net5),
    .A1(_3039_),
    .S(_1950_),
    .X(_1956_));
 sky130_fd_sc_hd__and2_1 _5182_ (.A(_1956_),
    .B(_1952_),
    .X(_1957_));
 sky130_fd_sc_hd__clkbuf_1 _5183_ (.A(_1957_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _5184_ (.A0(net4),
    .A1(_3044_),
    .S(_1950_),
    .X(_1958_));
 sky130_fd_sc_hd__and2_1 _5185_ (.A(_1958_),
    .B(_1952_),
    .X(_1959_));
 sky130_fd_sc_hd__clkbuf_1 _5186_ (.A(_1959_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _5187_ (.A0(net3),
    .A1(_0518_),
    .S(_1950_),
    .X(_1960_));
 sky130_fd_sc_hd__and2_1 _5188_ (.A(_1960_),
    .B(_1952_),
    .X(_1961_));
 sky130_fd_sc_hd__clkbuf_1 _5189_ (.A(_1961_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _5190_ (.A0(net2),
    .A1(_3037_),
    .S(_1950_),
    .X(_1962_));
 sky130_fd_sc_hd__and2_1 _5191_ (.A(_1962_),
    .B(_1952_),
    .X(_1963_));
 sky130_fd_sc_hd__clkbuf_1 _5192_ (.A(_1963_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(net16),
    .A1(_0516_),
    .S(_1950_),
    .X(_1964_));
 sky130_fd_sc_hd__and2_1 _5194_ (.A(_1964_),
    .B(_1952_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_1 _5195_ (.A(_1965_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _5196_ (.A0(net15),
    .A1(\BitStream_buffer.BS_buffer[7] ),
    .S(_1950_),
    .X(_1966_));
 sky130_fd_sc_hd__and2_1 _5197_ (.A(_1966_),
    .B(_1952_),
    .X(_1967_));
 sky130_fd_sc_hd__clkbuf_1 _5198_ (.A(_1967_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _5199_ (.A0(net14),
    .A1(_0330_),
    .S(_1950_),
    .X(_1968_));
 sky130_fd_sc_hd__and2_1 _5200_ (.A(_1968_),
    .B(_1952_),
    .X(_1969_));
 sky130_fd_sc_hd__clkbuf_1 _5201_ (.A(_1969_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(net13),
    .A1(_0325_),
    .S(_1950_),
    .X(_1970_));
 sky130_fd_sc_hd__and2_1 _5203_ (.A(_1970_),
    .B(_1952_),
    .X(_1971_));
 sky130_fd_sc_hd__clkbuf_1 _5204_ (.A(_1971_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _5205_ (.A0(net12),
    .A1(_0527_),
    .S(_1949_),
    .X(_1972_));
 sky130_fd_sc_hd__buf_2 _5206_ (.A(_0404_),
    .X(_1973_));
 sky130_fd_sc_hd__and2_1 _5207_ (.A(_1972_),
    .B(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__clkbuf_1 _5208_ (.A(_1974_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _5209_ (.A0(net11),
    .A1(_0650_),
    .S(_1949_),
    .X(_1975_));
 sky130_fd_sc_hd__and2_1 _5210_ (.A(_1975_),
    .B(_1973_),
    .X(_1976_));
 sky130_fd_sc_hd__clkbuf_1 _5211_ (.A(_1976_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _5212_ (.A0(net10),
    .A1(_0770_),
    .S(_1949_),
    .X(_1977_));
 sky130_fd_sc_hd__and2_1 _5213_ (.A(_1977_),
    .B(_1973_),
    .X(_1978_));
 sky130_fd_sc_hd__clkbuf_1 _5214_ (.A(_1978_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _5215_ (.A0(net9),
    .A1(_3051_),
    .S(_1949_),
    .X(_1979_));
 sky130_fd_sc_hd__and2_1 _5216_ (.A(_1979_),
    .B(_1973_),
    .X(_1980_));
 sky130_fd_sc_hd__clkbuf_1 _5217_ (.A(_1980_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _5218_ (.A0(net8),
    .A1(_0521_),
    .S(_1949_),
    .X(_1981_));
 sky130_fd_sc_hd__and2_1 _5219_ (.A(_1981_),
    .B(_1973_),
    .X(_1982_));
 sky130_fd_sc_hd__clkbuf_1 _5220_ (.A(_1982_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _5221_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[15] ),
    .S(_1949_),
    .X(_1983_));
 sky130_fd_sc_hd__and2_1 _5222_ (.A(_1983_),
    .B(_1973_),
    .X(_1984_));
 sky130_fd_sc_hd__clkbuf_1 _5223_ (.A(_1984_),
    .X(_0291_));
 sky130_fd_sc_hd__nor2_1 _5224_ (.A(net33),
    .B(_1936_),
    .Y(_1985_));
 sky130_fd_sc_hd__inv_2 _5225_ (.A(net31),
    .Y(_1986_));
 sky130_fd_sc_hd__and3_1 _5226_ (.A(_1985_),
    .B(net32),
    .C(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__o21ai_1 _5227_ (.A1(_0403_),
    .A2(_1987_),
    .B1(_0405_),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_2 _5228_ (.A(net29),
    .Y(_1988_));
 sky130_fd_sc_hd__nor2_1 _5229_ (.A(net28),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__nor2_1 _5230_ (.A(net28),
    .B(_1941_),
    .Y(_1990_));
 sky130_fd_sc_hd__and3_1 _5231_ (.A(_1946_),
    .B(_1947_),
    .C(\BitStream_buffer.buffer_index[6] ),
    .X(_1991_));
 sky130_fd_sc_hd__and4_1 _5232_ (.A(_3012_),
    .B(_2708_),
    .C(_1990_),
    .D(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__a31oi_2 _5233_ (.A1(\BitStream_buffer.pc[6] ),
    .A2(_1948_),
    .A3(_1990_),
    .B1(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__and4_1 _5234_ (.A(\BitStream_buffer.pc_previous[1] ),
    .B(\BitStream_buffer.pc_previous[0] ),
    .C(\BitStream_buffer.pc_previous[2] ),
    .D(\BitStream_buffer.pc_previous[3] ),
    .X(_1994_));
 sky130_fd_sc_hd__a31o_1 _5235_ (.A1(_1994_),
    .A2(\BitStream_buffer.pc_previous[4] ),
    .A3(\BitStream_buffer.pc_previous[5] ),
    .B1(\BitStream_buffer.pc_previous[6] ),
    .X(_1995_));
 sky130_fd_sc_hd__nor2_1 _5236_ (.A(\BitStream_buffer.pc_previous[6] ),
    .B(_2708_),
    .Y(_1996_));
 sky130_fd_sc_hd__a31o_1 _5237_ (.A1(_1995_),
    .A2(_2708_),
    .A3(_3012_),
    .B1(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__nand2_1 _5238_ (.A(_1997_),
    .B(_1990_),
    .Y(_1998_));
 sky130_fd_sc_hd__o21ai_1 _5239_ (.A1(net28),
    .A2(_1941_),
    .B1(_1942_),
    .Y(_1999_));
 sky130_fd_sc_hd__nand3_1 _5240_ (.A(_1993_),
    .B(_1998_),
    .C(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__nand2_2 _5241_ (.A(_2000_),
    .B(_1987_),
    .Y(_2001_));
 sky130_fd_sc_hd__a2111o_1 _5242_ (.A1(net30),
    .A2(net28),
    .B1(_1940_),
    .C1(_1989_),
    .D1(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_2001_),
    .B(net30),
    .Y(_2003_));
 sky130_fd_sc_hd__a21oi_1 _5244_ (.A1(_2002_),
    .A2(_2003_),
    .B1(_0675_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _5245_ (.A(_1988_),
    .B(net28),
    .Y(_2004_));
 sky130_fd_sc_hd__inv_2 _5246_ (.A(_1989_),
    .Y(_2005_));
 sky130_fd_sc_hd__a211o_1 _5247_ (.A1(_2004_),
    .A2(_2005_),
    .B1(net30),
    .C1(_2001_),
    .X(_2006_));
 sky130_fd_sc_hd__nand2_1 _5248_ (.A(_2001_),
    .B(net29),
    .Y(_2007_));
 sky130_fd_sc_hd__a21oi_1 _5249_ (.A1(_2006_),
    .A2(_2007_),
    .B1(_0675_),
    .Y(_0288_));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(net28),
    .B(_1943_),
    .X(_2008_));
 sky130_fd_sc_hd__a31o_1 _5251_ (.A1(_1998_),
    .A2(_1993_),
    .A3(_2008_),
    .B1(_2001_),
    .X(_2009_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(_2001_),
    .B(net28),
    .Y(_2010_));
 sky130_fd_sc_hd__a21oi_1 _5253_ (.A1(_2009_),
    .A2(_2010_),
    .B1(_0675_),
    .Y(_0287_));
 sky130_fd_sc_hd__nand2_1 _5254_ (.A(net32),
    .B(net31),
    .Y(_2011_));
 sky130_fd_sc_hd__inv_2 _5255_ (.A(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__a21o_1 _5256_ (.A1(_2012_),
    .A2(net33),
    .B1(net34),
    .X(_2013_));
 sky130_fd_sc_hd__inv_2 _5257_ (.A(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__nor2_1 _5258_ (.A(_0675_),
    .B(_2014_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_1 _5259_ (.A1(net33),
    .A2(_2012_),
    .B1(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__nand2_1 _5260_ (.A(net34),
    .B(net33),
    .Y(_2016_));
 sky130_fd_sc_hd__a21oi_1 _5261_ (.A1(_2015_),
    .A2(_2016_),
    .B1(_0675_),
    .Y(_0285_));
 sky130_fd_sc_hd__nor2_1 _5262_ (.A(_1986_),
    .B(_1938_),
    .Y(_2017_));
 sky130_fd_sc_hd__a21o_1 _5263_ (.A1(_2017_),
    .A2(net32),
    .B1(_0673_),
    .X(_2018_));
 sky130_fd_sc_hd__o21ba_1 _5264_ (.A1(net32),
    .A2(_2017_),
    .B1_N(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__clkbuf_1 _5265_ (.A(_2019_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _5266_ (.A(_0673_),
    .B(_2017_),
    .X(_2020_));
 sky130_fd_sc_hd__a21o_1 _5267_ (.A1(_1986_),
    .A2(_1938_),
    .B1(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__inv_2 _5268_ (.A(_2021_),
    .Y(_0283_));
 sky130_fd_sc_hd__or4b_1 _5269_ (.A(\BitStream_buffer.buffer_index[6] ),
    .B(_1946_),
    .C(\BitStream_buffer.buffer_index[4] ),
    .D_N(_1944_),
    .X(_2022_));
 sky130_fd_sc_hd__clkbuf_4 _5270_ (.A(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__clkbuf_4 _5271_ (.A(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(net7),
    .A1(\BitStream_buffer.BS_buffer[32] ),
    .S(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__and2_1 _5273_ (.A(_2025_),
    .B(_1973_),
    .X(_2026_));
 sky130_fd_sc_hd__clkbuf_1 _5274_ (.A(_2026_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5275_ (.A0(net6),
    .A1(\BitStream_buffer.BS_buffer[33] ),
    .S(_2024_),
    .X(_2027_));
 sky130_fd_sc_hd__and2_1 _5276_ (.A(_2027_),
    .B(_1973_),
    .X(_2028_));
 sky130_fd_sc_hd__clkbuf_1 _5277_ (.A(_2028_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(net5),
    .A1(\BitStream_buffer.BS_buffer[34] ),
    .S(_2024_),
    .X(_2029_));
 sky130_fd_sc_hd__and2_1 _5279_ (.A(_2029_),
    .B(_1973_),
    .X(_2030_));
 sky130_fd_sc_hd__clkbuf_1 _5280_ (.A(_2030_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(net4),
    .A1(\BitStream_buffer.BS_buffer[35] ),
    .S(_2024_),
    .X(_2031_));
 sky130_fd_sc_hd__and2_1 _5282_ (.A(_2031_),
    .B(_1973_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _5283_ (.A(_2032_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(net3),
    .A1(\BitStream_buffer.BS_buffer[36] ),
    .S(_2024_),
    .X(_2033_));
 sky130_fd_sc_hd__buf_2 _5285_ (.A(_0404_),
    .X(_2034_));
 sky130_fd_sc_hd__and2_1 _5286_ (.A(_2033_),
    .B(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _5287_ (.A(_2035_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5288_ (.A0(net2),
    .A1(\BitStream_buffer.BS_buffer[37] ),
    .S(_2024_),
    .X(_2036_));
 sky130_fd_sc_hd__and2_1 _5289_ (.A(_2036_),
    .B(_2034_),
    .X(_2037_));
 sky130_fd_sc_hd__clkbuf_1 _5290_ (.A(_2037_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(net16),
    .A1(\BitStream_buffer.BS_buffer[38] ),
    .S(_2024_),
    .X(_2038_));
 sky130_fd_sc_hd__and2_1 _5292_ (.A(_2038_),
    .B(_2034_),
    .X(_2039_));
 sky130_fd_sc_hd__clkbuf_1 _5293_ (.A(_2039_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(net15),
    .A1(\BitStream_buffer.BS_buffer[39] ),
    .S(_2024_),
    .X(_2040_));
 sky130_fd_sc_hd__and2_1 _5295_ (.A(_2040_),
    .B(_2034_),
    .X(_2041_));
 sky130_fd_sc_hd__clkbuf_1 _5296_ (.A(_2041_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(net14),
    .A1(\BitStream_buffer.BS_buffer[40] ),
    .S(_2024_),
    .X(_2042_));
 sky130_fd_sc_hd__and2_1 _5298_ (.A(_2042_),
    .B(_2034_),
    .X(_2043_));
 sky130_fd_sc_hd__clkbuf_1 _5299_ (.A(_2043_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(net13),
    .A1(\BitStream_buffer.BS_buffer[41] ),
    .S(_2024_),
    .X(_2044_));
 sky130_fd_sc_hd__and2_1 _5301_ (.A(_2044_),
    .B(_2034_),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_1 _5302_ (.A(_2045_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(net12),
    .A1(\BitStream_buffer.BS_buffer[42] ),
    .S(_2023_),
    .X(_2046_));
 sky130_fd_sc_hd__and2_1 _5304_ (.A(_2046_),
    .B(_2034_),
    .X(_2047_));
 sky130_fd_sc_hd__clkbuf_1 _5305_ (.A(_2047_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5306_ (.A0(net11),
    .A1(\BitStream_buffer.BS_buffer[43] ),
    .S(_2023_),
    .X(_2048_));
 sky130_fd_sc_hd__and2_1 _5307_ (.A(_2048_),
    .B(_2034_),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_1 _5308_ (.A(_2049_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net10),
    .A1(\BitStream_buffer.BS_buffer[44] ),
    .S(_2023_),
    .X(_2050_));
 sky130_fd_sc_hd__and2_1 _5310_ (.A(_2050_),
    .B(_2034_),
    .X(_2051_));
 sky130_fd_sc_hd__clkbuf_1 _5311_ (.A(_2051_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(net9),
    .A1(\BitStream_buffer.BS_buffer[45] ),
    .S(_2023_),
    .X(_2052_));
 sky130_fd_sc_hd__and2_1 _5313_ (.A(_2052_),
    .B(_2034_),
    .X(_2053_));
 sky130_fd_sc_hd__clkbuf_1 _5314_ (.A(_2053_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5315_ (.A0(net8),
    .A1(\BitStream_buffer.BS_buffer[46] ),
    .S(_2023_),
    .X(_2054_));
 sky130_fd_sc_hd__buf_2 _5316_ (.A(_0404_),
    .X(_2055_));
 sky130_fd_sc_hd__and2_1 _5317_ (.A(_2054_),
    .B(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__clkbuf_1 _5318_ (.A(_2056_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[47] ),
    .S(_2023_),
    .X(_2057_));
 sky130_fd_sc_hd__and2_1 _5320_ (.A(_2057_),
    .B(_2055_),
    .X(_2058_));
 sky130_fd_sc_hd__clkbuf_1 _5321_ (.A(_2058_),
    .X(_0267_));
 sky130_fd_sc_hd__or4b_1 _5322_ (.A(\BitStream_buffer.buffer_index[6] ),
    .B(\BitStream_buffer.buffer_index[5] ),
    .C(_1947_),
    .D_N(_1944_),
    .X(_2059_));
 sky130_fd_sc_hd__buf_2 _5323_ (.A(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__clkbuf_4 _5324_ (.A(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(net7),
    .A1(_0363_),
    .S(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__and2_1 _5326_ (.A(_2062_),
    .B(_2055_),
    .X(_2063_));
 sky130_fd_sc_hd__clkbuf_1 _5327_ (.A(_2063_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5328_ (.A0(net6),
    .A1(_0366_),
    .S(_2061_),
    .X(_2064_));
 sky130_fd_sc_hd__and2_1 _5329_ (.A(_2064_),
    .B(_2055_),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _5330_ (.A(_2065_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(net5),
    .A1(\BitStream_buffer.BS_buffer[18] ),
    .S(_2061_),
    .X(_2066_));
 sky130_fd_sc_hd__and2_1 _5332_ (.A(_2066_),
    .B(_2055_),
    .X(_2067_));
 sky130_fd_sc_hd__clkbuf_1 _5333_ (.A(_2067_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(net4),
    .A1(\BitStream_buffer.BS_buffer[19] ),
    .S(_2061_),
    .X(_2068_));
 sky130_fd_sc_hd__and2_1 _5335_ (.A(_2068_),
    .B(_2055_),
    .X(_2069_));
 sky130_fd_sc_hd__clkbuf_1 _5336_ (.A(_2069_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(net3),
    .A1(\BitStream_buffer.BS_buffer[20] ),
    .S(_2061_),
    .X(_2070_));
 sky130_fd_sc_hd__and2_1 _5338_ (.A(_2070_),
    .B(_2055_),
    .X(_2071_));
 sky130_fd_sc_hd__clkbuf_1 _5339_ (.A(_2071_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5340_ (.A0(net2),
    .A1(\BitStream_buffer.BS_buffer[21] ),
    .S(_2061_),
    .X(_2072_));
 sky130_fd_sc_hd__and2_1 _5341_ (.A(_2072_),
    .B(_2055_),
    .X(_2073_));
 sky130_fd_sc_hd__clkbuf_1 _5342_ (.A(_2073_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(net16),
    .A1(\BitStream_buffer.BS_buffer[22] ),
    .S(_2061_),
    .X(_2074_));
 sky130_fd_sc_hd__and2_1 _5344_ (.A(_2074_),
    .B(_2055_),
    .X(_2075_));
 sky130_fd_sc_hd__clkbuf_1 _5345_ (.A(_2075_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net15),
    .A1(\BitStream_buffer.BS_buffer[23] ),
    .S(_2061_),
    .X(_2076_));
 sky130_fd_sc_hd__and2_1 _5347_ (.A(_2076_),
    .B(_2055_),
    .X(_2077_));
 sky130_fd_sc_hd__clkbuf_1 _5348_ (.A(_2077_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5349_ (.A0(net14),
    .A1(\BitStream_buffer.BS_buffer[24] ),
    .S(_2061_),
    .X(_2078_));
 sky130_fd_sc_hd__buf_2 _5350_ (.A(_0404_),
    .X(_2079_));
 sky130_fd_sc_hd__and2_1 _5351_ (.A(_2078_),
    .B(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__clkbuf_1 _5352_ (.A(_2080_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(net13),
    .A1(\BitStream_buffer.BS_buffer[25] ),
    .S(_2061_),
    .X(_2081_));
 sky130_fd_sc_hd__and2_1 _5354_ (.A(_2081_),
    .B(_2079_),
    .X(_2082_));
 sky130_fd_sc_hd__clkbuf_1 _5355_ (.A(_2082_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(net12),
    .A1(\BitStream_buffer.BS_buffer[26] ),
    .S(_2060_),
    .X(_2083_));
 sky130_fd_sc_hd__and2_1 _5357_ (.A(_2083_),
    .B(_2079_),
    .X(_2084_));
 sky130_fd_sc_hd__clkbuf_1 _5358_ (.A(_2084_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5359_ (.A0(net11),
    .A1(\BitStream_buffer.BS_buffer[27] ),
    .S(_2060_),
    .X(_2085_));
 sky130_fd_sc_hd__and2_1 _5360_ (.A(_2085_),
    .B(_2079_),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_1 _5361_ (.A(_2086_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(net10),
    .A1(\BitStream_buffer.BS_buffer[28] ),
    .S(_2060_),
    .X(_2087_));
 sky130_fd_sc_hd__and2_1 _5363_ (.A(_2087_),
    .B(_2079_),
    .X(_2088_));
 sky130_fd_sc_hd__clkbuf_1 _5364_ (.A(_2088_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(net9),
    .A1(_0380_),
    .S(_2060_),
    .X(_2089_));
 sky130_fd_sc_hd__and2_1 _5366_ (.A(_2089_),
    .B(_2079_),
    .X(_2090_));
 sky130_fd_sc_hd__clkbuf_1 _5367_ (.A(_2090_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(net8),
    .A1(_0387_),
    .S(_2060_),
    .X(_2091_));
 sky130_fd_sc_hd__and2_1 _5369_ (.A(_2091_),
    .B(_2079_),
    .X(_2092_));
 sky130_fd_sc_hd__clkbuf_1 _5370_ (.A(_2092_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[31] ),
    .S(_2060_),
    .X(_2093_));
 sky130_fd_sc_hd__and2_1 _5372_ (.A(_2093_),
    .B(_2079_),
    .X(_2094_));
 sky130_fd_sc_hd__clkbuf_1 _5373_ (.A(_2094_),
    .X(_0251_));
 sky130_fd_sc_hd__or2_1 _5374_ (.A(\BitStream_buffer.pc_previous[1] ),
    .B(\BitStream_buffer.exp_golomb_len[1] ),
    .X(_2095_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(\BitStream_buffer.pc_previous[1] ),
    .B(\BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_2 _5376_ (.A(_2095_),
    .B(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__o21ai_4 _5377_ (.A1(_2611_),
    .A2(_2097_),
    .B1(_2096_),
    .Y(_2098_));
 sky130_fd_sc_hd__or2_1 _5378_ (.A(\BitStream_buffer.pc_previous[2] ),
    .B(\BitStream_buffer.exp_golomb_len[2] ),
    .X(_2099_));
 sky130_fd_sc_hd__nand2_1 _5379_ (.A(\BitStream_buffer.pc_previous[2] ),
    .B(\BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2100_));
 sky130_fd_sc_hd__a21bo_1 _5380_ (.A1(_2098_),
    .A2(_2099_),
    .B1_N(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__o21ai_1 _5381_ (.A1(\BitStream_buffer.pc_previous[3] ),
    .A2(\BitStream_buffer.exp_golomb_len[3] ),
    .B1(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand2_1 _5382_ (.A(\BitStream_buffer.pc_previous[3] ),
    .B(\BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2103_));
 sky130_fd_sc_hd__nand2_2 _5383_ (.A(_2102_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__and3_2 _5384_ (.A(_2104_),
    .B(\BitStream_buffer.pc_previous[4] ),
    .C(\BitStream_buffer.pc_previous[5] ),
    .X(_2105_));
 sky130_fd_sc_hd__xor2_4 _5385_ (.A(\BitStream_buffer.pc_previous[6] ),
    .B(_2105_),
    .X(\BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nand2_1 _5386_ (.A(_0405_),
    .B(\BitStream_buffer.pc[6] ),
    .Y(_2106_));
 sky130_fd_sc_hd__inv_2 _5387_ (.A(_2106_),
    .Y(_0250_));
 sky130_fd_sc_hd__a21oi_1 _5388_ (.A1(_2104_),
    .A2(\BitStream_buffer.pc_previous[4] ),
    .B1(\BitStream_buffer.pc_previous[5] ),
    .Y(_2107_));
 sky130_fd_sc_hd__nor2_2 _5389_ (.A(_2107_),
    .B(_2105_),
    .Y(\BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(_0405_),
    .B(\BitStream_buffer.pc[5] ),
    .Y(_2108_));
 sky130_fd_sc_hd__inv_2 _5391_ (.A(_2108_),
    .Y(_0249_));
 sky130_fd_sc_hd__xor2_4 _5392_ (.A(\BitStream_buffer.pc_previous[4] ),
    .B(_2104_),
    .X(\BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__nand2_1 _5393_ (.A(_0405_),
    .B(\BitStream_buffer.pc[4] ),
    .Y(_2109_));
 sky130_fd_sc_hd__inv_2 _5394_ (.A(_2109_),
    .Y(_0248_));
 sky130_fd_sc_hd__nor2_1 _5395_ (.A(\BitStream_buffer.pc_previous[3] ),
    .B(\BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2110_));
 sky130_fd_sc_hd__and2b_2 _5396_ (.A_N(_2110_),
    .B(_2103_),
    .X(_2111_));
 sky130_fd_sc_hd__xor2_4 _5397_ (.A(_2111_),
    .B(_2101_),
    .X(\BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__nand2_1 _5398_ (.A(_0405_),
    .B(\BitStream_buffer.pc[3] ),
    .Y(_2112_));
 sky130_fd_sc_hd__inv_2 _5399_ (.A(_2112_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_2 _5400_ (.A(_2099_),
    .B(_2100_),
    .Y(_2113_));
 sky130_fd_sc_hd__xnor2_4 _5401_ (.A(_2113_),
    .B(_2098_),
    .Y(\BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(_0405_),
    .B(\BitStream_buffer.pc[2] ),
    .Y(_2114_));
 sky130_fd_sc_hd__inv_2 _5403_ (.A(_2114_),
    .Y(_0246_));
 sky130_fd_sc_hd__xor2_4 _5404_ (.A(_2611_),
    .B(_2097_),
    .X(\BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__nand2_1 _5405_ (.A(_0405_),
    .B(\BitStream_buffer.pc[1] ),
    .Y(_2115_));
 sky130_fd_sc_hd__inv_2 _5406_ (.A(_2115_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand2_1 _5407_ (.A(_2618_),
    .B(_0405_),
    .Y(_2116_));
 sky130_fd_sc_hd__inv_2 _5408_ (.A(_2116_),
    .Y(_0244_));
 sky130_fd_sc_hd__nand2_1 _5409_ (.A(net201),
    .B(\BitStream_buffer.buffer_index[4] ),
    .Y(_2117_));
 sky130_fd_sc_hd__or2_1 _5410_ (.A(_1946_),
    .B(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__or2_1 _5411_ (.A(\BitStream_buffer.buffer_index[6] ),
    .B(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__clkbuf_4 _5412_ (.A(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__buf_4 _5413_ (.A(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__mux2_1 _5414_ (.A0(net7),
    .A1(\BitStream_buffer.BS_buffer[48] ),
    .S(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__and2_1 _5415_ (.A(_2122_),
    .B(_2079_),
    .X(_2123_));
 sky130_fd_sc_hd__clkbuf_1 _5416_ (.A(_2123_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5417_ (.A0(net6),
    .A1(\BitStream_buffer.BS_buffer[49] ),
    .S(_2121_),
    .X(_2124_));
 sky130_fd_sc_hd__and2_1 _5418_ (.A(_2124_),
    .B(_2079_),
    .X(_2125_));
 sky130_fd_sc_hd__clkbuf_1 _5419_ (.A(_2125_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5420_ (.A0(net5),
    .A1(\BitStream_buffer.BS_buffer[50] ),
    .S(_2121_),
    .X(_2126_));
 sky130_fd_sc_hd__clkbuf_2 _5421_ (.A(_0404_),
    .X(_2127_));
 sky130_fd_sc_hd__and2_1 _5422_ (.A(_2126_),
    .B(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _5423_ (.A(_2128_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(net4),
    .A1(\BitStream_buffer.BS_buffer[51] ),
    .S(_2121_),
    .X(_2129_));
 sky130_fd_sc_hd__and2_1 _5425_ (.A(_2129_),
    .B(_2127_),
    .X(_2130_));
 sky130_fd_sc_hd__clkbuf_1 _5426_ (.A(_2130_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5427_ (.A0(net3),
    .A1(\BitStream_buffer.BS_buffer[52] ),
    .S(_2121_),
    .X(_2131_));
 sky130_fd_sc_hd__and2_1 _5428_ (.A(_2131_),
    .B(_2127_),
    .X(_2132_));
 sky130_fd_sc_hd__clkbuf_1 _5429_ (.A(_2132_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5430_ (.A0(net2),
    .A1(\BitStream_buffer.BS_buffer[53] ),
    .S(_2121_),
    .X(_2133_));
 sky130_fd_sc_hd__and2_1 _5431_ (.A(_2133_),
    .B(_2127_),
    .X(_2134_));
 sky130_fd_sc_hd__clkbuf_1 _5432_ (.A(_2134_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(net16),
    .A1(\BitStream_buffer.BS_buffer[54] ),
    .S(_2121_),
    .X(_2135_));
 sky130_fd_sc_hd__and2_1 _5434_ (.A(_2135_),
    .B(_2127_),
    .X(_2136_));
 sky130_fd_sc_hd__clkbuf_1 _5435_ (.A(_2136_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(net15),
    .A1(\BitStream_buffer.BS_buffer[55] ),
    .S(_2121_),
    .X(_2137_));
 sky130_fd_sc_hd__and2_1 _5437_ (.A(_2137_),
    .B(_2127_),
    .X(_2138_));
 sky130_fd_sc_hd__clkbuf_1 _5438_ (.A(_2138_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5439_ (.A0(net14),
    .A1(\BitStream_buffer.BS_buffer[56] ),
    .S(_2121_),
    .X(_2139_));
 sky130_fd_sc_hd__and2_1 _5440_ (.A(_2139_),
    .B(_2127_),
    .X(_2140_));
 sky130_fd_sc_hd__clkbuf_1 _5441_ (.A(_2140_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(net13),
    .A1(\BitStream_buffer.BS_buffer[57] ),
    .S(_2120_),
    .X(_2141_));
 sky130_fd_sc_hd__and2_1 _5443_ (.A(_2141_),
    .B(_2127_),
    .X(_2142_));
 sky130_fd_sc_hd__clkbuf_1 _5444_ (.A(_2142_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5445_ (.A0(net12),
    .A1(\BitStream_buffer.BS_buffer[58] ),
    .S(_2120_),
    .X(_2143_));
 sky130_fd_sc_hd__and2_1 _5446_ (.A(_2143_),
    .B(_2127_),
    .X(_2144_));
 sky130_fd_sc_hd__clkbuf_1 _5447_ (.A(_2144_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5448_ (.A0(net11),
    .A1(\BitStream_buffer.BS_buffer[59] ),
    .S(_2120_),
    .X(_2145_));
 sky130_fd_sc_hd__and2_1 _5449_ (.A(_2145_),
    .B(_2127_),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_1 _5450_ (.A(_2146_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5451_ (.A0(net10),
    .A1(\BitStream_buffer.BS_buffer[60] ),
    .S(_2120_),
    .X(_2147_));
 sky130_fd_sc_hd__clkbuf_2 _5452_ (.A(_0404_),
    .X(_2148_));
 sky130_fd_sc_hd__and2_1 _5453_ (.A(_2147_),
    .B(_2148_),
    .X(_2149_));
 sky130_fd_sc_hd__clkbuf_1 _5454_ (.A(_2149_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(net9),
    .A1(\BitStream_buffer.BS_buffer[61] ),
    .S(_2120_),
    .X(_2150_));
 sky130_fd_sc_hd__and2_1 _5456_ (.A(_2150_),
    .B(_2148_),
    .X(_2151_));
 sky130_fd_sc_hd__clkbuf_1 _5457_ (.A(_2151_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5458_ (.A0(net8),
    .A1(\BitStream_buffer.BS_buffer[62] ),
    .S(_2120_),
    .X(_2152_));
 sky130_fd_sc_hd__and2_1 _5459_ (.A(_2152_),
    .B(_2148_),
    .X(_2153_));
 sky130_fd_sc_hd__clkbuf_1 _5460_ (.A(_2153_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[63] ),
    .S(_2120_),
    .X(_2154_));
 sky130_fd_sc_hd__and2_1 _5462_ (.A(_2154_),
    .B(_2148_),
    .X(_2155_));
 sky130_fd_sc_hd__clkbuf_1 _5463_ (.A(_2155_),
    .X(_0228_));
 sky130_fd_sc_hd__nand2_4 _5464_ (.A(_1944_),
    .B(_1991_),
    .Y(_2156_));
 sky130_fd_sc_hd__clkbuf_4 _5465_ (.A(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__mux2_1 _5466_ (.A0(net7),
    .A1(\BitStream_buffer.BS_buffer[64] ),
    .S(_2157_),
    .X(_2158_));
 sky130_fd_sc_hd__and2_1 _5467_ (.A(_2158_),
    .B(_2148_),
    .X(_2159_));
 sky130_fd_sc_hd__clkbuf_1 _5468_ (.A(_2159_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(net6),
    .A1(\BitStream_buffer.BS_buffer[65] ),
    .S(_2157_),
    .X(_2160_));
 sky130_fd_sc_hd__and2_1 _5470_ (.A(_2160_),
    .B(_2148_),
    .X(_2161_));
 sky130_fd_sc_hd__clkbuf_1 _5471_ (.A(_2161_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(net5),
    .A1(\BitStream_buffer.BS_buffer[66] ),
    .S(_2157_),
    .X(_2162_));
 sky130_fd_sc_hd__and2_1 _5473_ (.A(_2162_),
    .B(_2148_),
    .X(_2163_));
 sky130_fd_sc_hd__clkbuf_1 _5474_ (.A(_2163_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5475_ (.A0(net4),
    .A1(\BitStream_buffer.BS_buffer[67] ),
    .S(_2157_),
    .X(_2164_));
 sky130_fd_sc_hd__and2_1 _5476_ (.A(_2164_),
    .B(_2148_),
    .X(_2165_));
 sky130_fd_sc_hd__clkbuf_1 _5477_ (.A(_2165_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(net3),
    .A1(\BitStream_buffer.BS_buffer[68] ),
    .S(_2157_),
    .X(_2166_));
 sky130_fd_sc_hd__and2_1 _5479_ (.A(_2166_),
    .B(_2148_),
    .X(_2167_));
 sky130_fd_sc_hd__clkbuf_1 _5480_ (.A(_2167_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5481_ (.A0(net2),
    .A1(\BitStream_buffer.BS_buffer[69] ),
    .S(_2157_),
    .X(_2168_));
 sky130_fd_sc_hd__and2_1 _5482_ (.A(_2168_),
    .B(_2148_),
    .X(_2169_));
 sky130_fd_sc_hd__clkbuf_1 _5483_ (.A(_2169_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(net16),
    .A1(\BitStream_buffer.BS_buffer[70] ),
    .S(_2157_),
    .X(_2170_));
 sky130_fd_sc_hd__buf_2 _5485_ (.A(_0404_),
    .X(_2171_));
 sky130_fd_sc_hd__and2_1 _5486_ (.A(_2170_),
    .B(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__clkbuf_1 _5487_ (.A(_2172_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(net15),
    .A1(\BitStream_buffer.BS_buffer[71] ),
    .S(_2157_),
    .X(_2173_));
 sky130_fd_sc_hd__and2_1 _5489_ (.A(_2173_),
    .B(_2171_),
    .X(_2174_));
 sky130_fd_sc_hd__clkbuf_1 _5490_ (.A(_2174_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5491_ (.A0(net14),
    .A1(\BitStream_buffer.BS_buffer[72] ),
    .S(_2157_),
    .X(_2175_));
 sky130_fd_sc_hd__and2_1 _5492_ (.A(_2175_),
    .B(_2171_),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_1 _5493_ (.A(_2176_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(net13),
    .A1(\BitStream_buffer.BS_buffer[73] ),
    .S(_2157_),
    .X(_2177_));
 sky130_fd_sc_hd__and2_1 _5495_ (.A(_2177_),
    .B(_2171_),
    .X(_2178_));
 sky130_fd_sc_hd__clkbuf_1 _5496_ (.A(_2178_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _5497_ (.A0(net12),
    .A1(\BitStream_buffer.BS_buffer[74] ),
    .S(_2156_),
    .X(_2179_));
 sky130_fd_sc_hd__and2_1 _5498_ (.A(_2179_),
    .B(_2171_),
    .X(_2180_));
 sky130_fd_sc_hd__clkbuf_1 _5499_ (.A(_2180_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(net11),
    .A1(\BitStream_buffer.BS_buffer[75] ),
    .S(_2156_),
    .X(_2181_));
 sky130_fd_sc_hd__and2_1 _5501_ (.A(_2181_),
    .B(_2171_),
    .X(_2182_));
 sky130_fd_sc_hd__clkbuf_1 _5502_ (.A(_2182_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5503_ (.A0(net10),
    .A1(\BitStream_buffer.BS_buffer[76] ),
    .S(_2156_),
    .X(_2183_));
 sky130_fd_sc_hd__and2_1 _5504_ (.A(_2183_),
    .B(_2171_),
    .X(_2184_));
 sky130_fd_sc_hd__clkbuf_1 _5505_ (.A(_2184_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5506_ (.A0(net9),
    .A1(\BitStream_buffer.BS_buffer[77] ),
    .S(_2156_),
    .X(_2185_));
 sky130_fd_sc_hd__and2_1 _5507_ (.A(_2185_),
    .B(_2171_),
    .X(_2186_));
 sky130_fd_sc_hd__clkbuf_1 _5508_ (.A(_2186_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(net8),
    .A1(\BitStream_buffer.BS_buffer[78] ),
    .S(_2156_),
    .X(_2187_));
 sky130_fd_sc_hd__and2_1 _5510_ (.A(_2187_),
    .B(_2171_),
    .X(_2188_));
 sky130_fd_sc_hd__clkbuf_1 _5511_ (.A(_2188_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[79] ),
    .S(_2156_),
    .X(_2189_));
 sky130_fd_sc_hd__and2_1 _5513_ (.A(_2189_),
    .B(_2171_),
    .X(_2190_));
 sky130_fd_sc_hd__clkbuf_1 _5514_ (.A(_2190_),
    .X(_0212_));
 sky130_fd_sc_hd__or4b_2 _5515_ (.A(_1945_),
    .B(\BitStream_buffer.buffer_index[5] ),
    .C(_1947_),
    .D_N(_1944_),
    .X(_2191_));
 sky130_fd_sc_hd__buf_2 _5516_ (.A(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__clkbuf_4 _5517_ (.A(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(net7),
    .A1(\BitStream_buffer.BS_buffer[80] ),
    .S(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__clkbuf_2 _5519_ (.A(_0404_),
    .X(_2195_));
 sky130_fd_sc_hd__and2_1 _5520_ (.A(_2194_),
    .B(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__clkbuf_1 _5521_ (.A(_2196_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(net6),
    .A1(\BitStream_buffer.BS_buffer[81] ),
    .S(_2193_),
    .X(_2197_));
 sky130_fd_sc_hd__and2_1 _5523_ (.A(_2197_),
    .B(_2195_),
    .X(_2198_));
 sky130_fd_sc_hd__clkbuf_1 _5524_ (.A(_2198_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _5525_ (.A0(net5),
    .A1(\BitStream_buffer.BS_buffer[82] ),
    .S(_2193_),
    .X(_2199_));
 sky130_fd_sc_hd__and2_1 _5526_ (.A(_2199_),
    .B(_2195_),
    .X(_2200_));
 sky130_fd_sc_hd__clkbuf_1 _5527_ (.A(_2200_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _5528_ (.A0(net4),
    .A1(\BitStream_buffer.BS_buffer[83] ),
    .S(_2193_),
    .X(_2201_));
 sky130_fd_sc_hd__and2_1 _5529_ (.A(_2201_),
    .B(_2195_),
    .X(_2202_));
 sky130_fd_sc_hd__clkbuf_1 _5530_ (.A(_2202_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _5531_ (.A0(net3),
    .A1(_2766_),
    .S(_2193_),
    .X(_2203_));
 sky130_fd_sc_hd__and2_1 _5532_ (.A(_2203_),
    .B(_2195_),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_1 _5533_ (.A(_2204_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(net2),
    .A1(_2768_),
    .S(_2193_),
    .X(_2205_));
 sky130_fd_sc_hd__and2_1 _5535_ (.A(_2205_),
    .B(_2195_),
    .X(_2206_));
 sky130_fd_sc_hd__clkbuf_1 _5536_ (.A(_2206_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _5537_ (.A0(net16),
    .A1(_2762_),
    .S(_2193_),
    .X(_2207_));
 sky130_fd_sc_hd__and2_1 _5538_ (.A(_2207_),
    .B(_2195_),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_1 _5539_ (.A(_2208_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _5540_ (.A0(net15),
    .A1(_2756_),
    .S(_2193_),
    .X(_2209_));
 sky130_fd_sc_hd__and2_1 _5541_ (.A(_2209_),
    .B(_2195_),
    .X(_2210_));
 sky130_fd_sc_hd__clkbuf_1 _5542_ (.A(_2210_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(net14),
    .A1(_2725_),
    .S(_2193_),
    .X(_2211_));
 sky130_fd_sc_hd__and2_1 _5544_ (.A(_2211_),
    .B(_2195_),
    .X(_2212_));
 sky130_fd_sc_hd__clkbuf_1 _5545_ (.A(_2212_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _5546_ (.A0(net13),
    .A1(_2706_),
    .S(_2193_),
    .X(_2213_));
 sky130_fd_sc_hd__and2_1 _5547_ (.A(_2213_),
    .B(_2195_),
    .X(_2214_));
 sky130_fd_sc_hd__clkbuf_1 _5548_ (.A(_2214_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _5549_ (.A0(net12),
    .A1(_2721_),
    .S(_2192_),
    .X(_2215_));
 sky130_fd_sc_hd__clkbuf_2 _5550_ (.A(net19),
    .X(_2216_));
 sky130_fd_sc_hd__and2_1 _5551_ (.A(_2215_),
    .B(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__clkbuf_1 _5552_ (.A(_2217_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _5553_ (.A0(net11),
    .A1(_2714_),
    .S(_2192_),
    .X(_2218_));
 sky130_fd_sc_hd__and2_1 _5554_ (.A(_2218_),
    .B(_2216_),
    .X(_2219_));
 sky130_fd_sc_hd__clkbuf_1 _5555_ (.A(_2219_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(net10),
    .A1(_2736_),
    .S(_2192_),
    .X(_2220_));
 sky130_fd_sc_hd__and2_1 _5557_ (.A(_2220_),
    .B(_2216_),
    .X(_2221_));
 sky130_fd_sc_hd__clkbuf_1 _5558_ (.A(_2221_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(net9),
    .A1(\BitStream_buffer.BS_buffer[93] ),
    .S(_2192_),
    .X(_2222_));
 sky130_fd_sc_hd__and2_1 _5560_ (.A(_2222_),
    .B(_2216_),
    .X(_2223_));
 sky130_fd_sc_hd__clkbuf_1 _5561_ (.A(_2223_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _5562_ (.A0(net8),
    .A1(\BitStream_buffer.BS_buffer[94] ),
    .S(_2192_),
    .X(_2224_));
 sky130_fd_sc_hd__and2_1 _5563_ (.A(_2224_),
    .B(_2216_),
    .X(_2225_));
 sky130_fd_sc_hd__clkbuf_1 _5564_ (.A(_2225_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[95] ),
    .S(_2192_),
    .X(_2226_));
 sky130_fd_sc_hd__and2_1 _5566_ (.A(_2226_),
    .B(_2216_),
    .X(_2227_));
 sky130_fd_sc_hd__clkbuf_1 _5567_ (.A(_2227_),
    .X(_0196_));
 sky130_fd_sc_hd__or4b_2 _5568_ (.A(_1945_),
    .B(_1946_),
    .C(\BitStream_buffer.buffer_index[4] ),
    .D_N(_1944_),
    .X(_2228_));
 sky130_fd_sc_hd__clkbuf_4 _5569_ (.A(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__clkbuf_4 _5570_ (.A(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(net7),
    .A1(_2800_),
    .S(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__and2_1 _5572_ (.A(_2231_),
    .B(_2216_),
    .X(_2232_));
 sky130_fd_sc_hd__clkbuf_1 _5573_ (.A(_2232_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(net6),
    .A1(\BitStream_buffer.BS_buffer[97] ),
    .S(_2230_),
    .X(_2233_));
 sky130_fd_sc_hd__and2_1 _5575_ (.A(_2233_),
    .B(_2216_),
    .X(_2234_));
 sky130_fd_sc_hd__clkbuf_1 _5576_ (.A(_2234_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _5577_ (.A0(net5),
    .A1(_2804_),
    .S(_2230_),
    .X(_2235_));
 sky130_fd_sc_hd__and2_1 _5578_ (.A(_2235_),
    .B(_2216_),
    .X(_2236_));
 sky130_fd_sc_hd__clkbuf_1 _5579_ (.A(_2236_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(net4),
    .A1(\BitStream_buffer.BS_buffer[99] ),
    .S(_2230_),
    .X(_2237_));
 sky130_fd_sc_hd__and2_1 _5581_ (.A(_2237_),
    .B(_2216_),
    .X(_2238_));
 sky130_fd_sc_hd__clkbuf_1 _5582_ (.A(_2238_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(net3),
    .A1(_2820_),
    .S(_2230_),
    .X(_2239_));
 sky130_fd_sc_hd__clkbuf_2 _5584_ (.A(net19),
    .X(_2240_));
 sky130_fd_sc_hd__and2_1 _5585_ (.A(_2239_),
    .B(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__clkbuf_1 _5586_ (.A(_2241_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(net2),
    .A1(\BitStream_buffer.BS_buffer[101] ),
    .S(_2230_),
    .X(_2242_));
 sky130_fd_sc_hd__and2_1 _5588_ (.A(_2242_),
    .B(_2240_),
    .X(_2243_));
 sky130_fd_sc_hd__clkbuf_1 _5589_ (.A(_2243_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _5590_ (.A0(net16),
    .A1(_2816_),
    .S(_2230_),
    .X(_2244_));
 sky130_fd_sc_hd__and2_1 _5591_ (.A(_2244_),
    .B(_2240_),
    .X(_2245_));
 sky130_fd_sc_hd__clkbuf_1 _5592_ (.A(_2245_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(net15),
    .A1(\BitStream_buffer.BS_buffer[103] ),
    .S(_2230_),
    .X(_2246_));
 sky130_fd_sc_hd__and2_1 _5594_ (.A(_2246_),
    .B(_2240_),
    .X(_2247_));
 sky130_fd_sc_hd__clkbuf_1 _5595_ (.A(_2247_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _5596_ (.A0(net14),
    .A1(_2792_),
    .S(_2230_),
    .X(_2248_));
 sky130_fd_sc_hd__and2_1 _5597_ (.A(_2248_),
    .B(_2240_),
    .X(_2249_));
 sky130_fd_sc_hd__clkbuf_1 _5598_ (.A(_2249_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(net13),
    .A1(\BitStream_buffer.BS_buffer[105] ),
    .S(_2230_),
    .X(_2250_));
 sky130_fd_sc_hd__and2_1 _5600_ (.A(_2250_),
    .B(_2240_),
    .X(_2251_));
 sky130_fd_sc_hd__clkbuf_1 _5601_ (.A(_2251_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _5602_ (.A0(net12),
    .A1(_2788_),
    .S(_2229_),
    .X(_2252_));
 sky130_fd_sc_hd__and2_1 _5603_ (.A(_2252_),
    .B(_2240_),
    .X(_2253_));
 sky130_fd_sc_hd__clkbuf_1 _5604_ (.A(_2253_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _5605_ (.A0(net11),
    .A1(_2781_),
    .S(_2229_),
    .X(_2254_));
 sky130_fd_sc_hd__and2_1 _5606_ (.A(_2254_),
    .B(_2240_),
    .X(_2255_));
 sky130_fd_sc_hd__clkbuf_1 _5607_ (.A(_2255_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _5608_ (.A0(net10),
    .A1(_2832_),
    .S(_2229_),
    .X(_2256_));
 sky130_fd_sc_hd__and2_1 _5609_ (.A(_2256_),
    .B(_2240_),
    .X(_2257_));
 sky130_fd_sc_hd__clkbuf_1 _5610_ (.A(_2257_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(net9),
    .A1(_2838_),
    .S(_2229_),
    .X(_2258_));
 sky130_fd_sc_hd__and2_1 _5612_ (.A(_2258_),
    .B(_2240_),
    .X(_2259_));
 sky130_fd_sc_hd__clkbuf_1 _5613_ (.A(_2259_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(net8),
    .A1(_2836_),
    .S(_2229_),
    .X(_2260_));
 sky130_fd_sc_hd__clkbuf_2 _5615_ (.A(net19),
    .X(_2261_));
 sky130_fd_sc_hd__and2_1 _5616_ (.A(_2260_),
    .B(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_1 _5617_ (.A(_2262_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _5618_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[111] ),
    .S(_2229_),
    .X(_2263_));
 sky130_fd_sc_hd__and2_1 _5619_ (.A(_2263_),
    .B(_2261_),
    .X(_2264_));
 sky130_fd_sc_hd__clkbuf_1 _5620_ (.A(_2264_),
    .X(_0180_));
 sky130_fd_sc_hd__or2_1 _5621_ (.A(_1945_),
    .B(_2118_),
    .X(_2265_));
 sky130_fd_sc_hd__buf_2 _5622_ (.A(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__clkbuf_4 _5623_ (.A(_2266_),
    .X(_2267_));
 sky130_fd_sc_hd__mux2_1 _5624_ (.A0(net7),
    .A1(\BitStream_buffer.BS_buffer[112] ),
    .S(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__and2_1 _5625_ (.A(_2268_),
    .B(_2261_),
    .X(_2269_));
 sky130_fd_sc_hd__clkbuf_1 _5626_ (.A(_2269_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _5627_ (.A0(net6),
    .A1(\BitStream_buffer.BS_buffer[113] ),
    .S(_2267_),
    .X(_2270_));
 sky130_fd_sc_hd__and2_1 _5628_ (.A(_2270_),
    .B(_2261_),
    .X(_2271_));
 sky130_fd_sc_hd__clkbuf_1 _5629_ (.A(_2271_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _5630_ (.A0(net5),
    .A1(\BitStream_buffer.BS_buffer[114] ),
    .S(_2267_),
    .X(_2272_));
 sky130_fd_sc_hd__and2_1 _5631_ (.A(_2272_),
    .B(_2261_),
    .X(_2273_));
 sky130_fd_sc_hd__clkbuf_1 _5632_ (.A(_2273_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _5633_ (.A0(net4),
    .A1(\BitStream_buffer.BS_buffer[115] ),
    .S(_2267_),
    .X(_2274_));
 sky130_fd_sc_hd__and2_1 _5634_ (.A(_2274_),
    .B(_2261_),
    .X(_2275_));
 sky130_fd_sc_hd__clkbuf_1 _5635_ (.A(_2275_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(net3),
    .A1(\BitStream_buffer.BS_buffer[116] ),
    .S(_2267_),
    .X(_2276_));
 sky130_fd_sc_hd__and2_1 _5637_ (.A(_2276_),
    .B(_2261_),
    .X(_2277_));
 sky130_fd_sc_hd__clkbuf_1 _5638_ (.A(_2277_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _5639_ (.A0(net2),
    .A1(\BitStream_buffer.BS_buffer[117] ),
    .S(_2267_),
    .X(_2278_));
 sky130_fd_sc_hd__and2_1 _5640_ (.A(_2278_),
    .B(_2261_),
    .X(_2279_));
 sky130_fd_sc_hd__clkbuf_1 _5641_ (.A(_2279_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5642_ (.A0(net16),
    .A1(\BitStream_buffer.BS_buffer[118] ),
    .S(_2267_),
    .X(_2280_));
 sky130_fd_sc_hd__and2_1 _5643_ (.A(_2280_),
    .B(_2261_),
    .X(_2281_));
 sky130_fd_sc_hd__clkbuf_1 _5644_ (.A(_2281_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _5645_ (.A0(net15),
    .A1(\BitStream_buffer.BS_buffer[119] ),
    .S(_2267_),
    .X(_2282_));
 sky130_fd_sc_hd__and2_1 _5646_ (.A(_2282_),
    .B(_2261_),
    .X(_2283_));
 sky130_fd_sc_hd__clkbuf_1 _5647_ (.A(_2283_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5648_ (.A0(net14),
    .A1(\BitStream_buffer.BS_buffer[120] ),
    .S(_2267_),
    .X(_2284_));
 sky130_fd_sc_hd__buf_2 _5649_ (.A(net19),
    .X(_2285_));
 sky130_fd_sc_hd__and2_1 _5650_ (.A(_2284_),
    .B(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__clkbuf_1 _5651_ (.A(_2286_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5652_ (.A0(net13),
    .A1(\BitStream_buffer.BS_buffer[121] ),
    .S(_2267_),
    .X(_2287_));
 sky130_fd_sc_hd__and2_1 _5653_ (.A(_2287_),
    .B(_2285_),
    .X(_2288_));
 sky130_fd_sc_hd__clkbuf_1 _5654_ (.A(_2288_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5655_ (.A0(net12),
    .A1(\BitStream_buffer.BS_buffer[122] ),
    .S(_2266_),
    .X(_2289_));
 sky130_fd_sc_hd__and2_1 _5656_ (.A(_2289_),
    .B(_2285_),
    .X(_2290_));
 sky130_fd_sc_hd__clkbuf_1 _5657_ (.A(_2290_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5658_ (.A0(net11),
    .A1(\BitStream_buffer.BS_buffer[123] ),
    .S(_2266_),
    .X(_2291_));
 sky130_fd_sc_hd__and2_1 _5659_ (.A(_2291_),
    .B(_2285_),
    .X(_2292_));
 sky130_fd_sc_hd__clkbuf_1 _5660_ (.A(_2292_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5661_ (.A0(net10),
    .A1(\BitStream_buffer.BS_buffer[124] ),
    .S(_2266_),
    .X(_2293_));
 sky130_fd_sc_hd__and2_1 _5662_ (.A(_2293_),
    .B(_2285_),
    .X(_2294_));
 sky130_fd_sc_hd__clkbuf_1 _5663_ (.A(_2294_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5664_ (.A0(net9),
    .A1(\BitStream_buffer.BS_buffer[125] ),
    .S(_2266_),
    .X(_2295_));
 sky130_fd_sc_hd__and2_1 _5665_ (.A(_2295_),
    .B(_2285_),
    .X(_2296_));
 sky130_fd_sc_hd__clkbuf_1 _5666_ (.A(_2296_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5667_ (.A0(net8),
    .A1(\BitStream_buffer.BS_buffer[126] ),
    .S(_2266_),
    .X(_2297_));
 sky130_fd_sc_hd__and2_1 _5668_ (.A(_2297_),
    .B(_2285_),
    .X(_2298_));
 sky130_fd_sc_hd__clkbuf_1 _5669_ (.A(_2298_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5670_ (.A0(net1),
    .A1(\BitStream_buffer.BS_buffer[127] ),
    .S(_2266_),
    .X(_2299_));
 sky130_fd_sc_hd__and2_1 _5671_ (.A(_2299_),
    .B(_2285_),
    .X(_2300_));
 sky130_fd_sc_hd__clkbuf_1 _5672_ (.A(_2300_),
    .X(_0164_));
 sky130_fd_sc_hd__nand2_1 _5673_ (.A(_2118_),
    .B(\BitStream_buffer.buffer_index[6] ),
    .Y(_2301_));
 sky130_fd_sc_hd__a21oi_1 _5674_ (.A1(_2121_),
    .A2(_2301_),
    .B1(_0675_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_2117_),
    .B(_1946_),
    .Y(_2302_));
 sky130_fd_sc_hd__and3_1 _5676_ (.A(_2118_),
    .B(_2285_),
    .C(_2302_),
    .X(_2303_));
 sky130_fd_sc_hd__clkbuf_1 _5677_ (.A(_2303_),
    .X(_0162_));
 sky130_fd_sc_hd__or2_1 _5678_ (.A(\BitStream_buffer.buffer_index[4] ),
    .B(_1944_),
    .X(_2304_));
 sky130_fd_sc_hd__and3_1 _5679_ (.A(_2304_),
    .B(_2285_),
    .C(_2117_),
    .X(_2305_));
 sky130_fd_sc_hd__clkbuf_1 _5680_ (.A(_2305_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _5681_ (.A(net18),
    .B(net17),
    .Y(_2306_));
 sky130_fd_sc_hd__inv_2 _5682_ (.A(_2306_),
    .Y(_2307_));
 sky130_fd_sc_hd__and3b_1 _5683_ (.A_N(net21),
    .B(_2307_),
    .C(net20),
    .X(_2308_));
 sky130_fd_sc_hd__inv_2 _5684_ (.A(\exp_golomb_decoding.te_range[2] ),
    .Y(_2309_));
 sky130_fd_sc_hd__and2_2 _5685_ (.A(_2308_),
    .B(_2309_),
    .X(_2310_));
 sky130_fd_sc_hd__nor2_1 _5686_ (.A(\BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2311_));
 sky130_fd_sc_hd__nand2_1 _5687_ (.A(_2311_),
    .B(_0403_),
    .Y(_2312_));
 sky130_fd_sc_hd__nand2_1 _5688_ (.A(_0787_),
    .B(_0894_),
    .Y(_2313_));
 sky130_fd_sc_hd__nor2_1 _5689_ (.A(\BitStream_buffer.BitStream_buffer_output[13] ),
    .B(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_2314_),
    .B(_0998_),
    .Y(_2315_));
 sky130_fd_sc_hd__inv_2 _5691_ (.A(_2315_),
    .Y(_2316_));
 sky130_fd_sc_hd__and3_1 _5692_ (.A(_2316_),
    .B(_1102_),
    .C(_1206_),
    .X(_2317_));
 sky130_fd_sc_hd__inv_2 _5693_ (.A(_2317_),
    .Y(_2318_));
 sky130_fd_sc_hd__nor2_1 _5694_ (.A(_2312_),
    .B(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__nor2_1 _5695_ (.A(\BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2320_));
 sky130_fd_sc_hd__inv_2 _5696_ (.A(_2320_),
    .Y(_2321_));
 sky130_fd_sc_hd__nor2_1 _5697_ (.A(\BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__nand2_1 _5698_ (.A(_2322_),
    .B(_1622_),
    .Y(_2323_));
 sky130_fd_sc_hd__inv_2 _5699_ (.A(_2312_),
    .Y(_2324_));
 sky130_fd_sc_hd__nor2_1 _5700_ (.A(\BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2325_));
 sky130_fd_sc_hd__nand2_2 _5701_ (.A(_2324_),
    .B(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__a21o_1 _5702_ (.A1(_2317_),
    .A2(_2323_),
    .B1(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__nor2_2 _5703_ (.A(_2319_),
    .B(_2327_),
    .Y(_2328_));
 sky130_fd_sc_hd__inv_6 _5704_ (.A(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__nand2_1 _5705_ (.A(_1830_),
    .B(\BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2330_));
 sky130_fd_sc_hd__nand2_1 _5706_ (.A(_2330_),
    .B(_1726_),
    .Y(_2331_));
 sky130_fd_sc_hd__nand2_1 _5707_ (.A(_2331_),
    .B(_1622_),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _5708_ (.A(_2332_),
    .B(_1518_),
    .Y(_2333_));
 sky130_fd_sc_hd__nand2_1 _5709_ (.A(_2333_),
    .B(_1414_),
    .Y(_2334_));
 sky130_fd_sc_hd__nand2_1 _5710_ (.A(_2334_),
    .B(_1310_),
    .Y(_2335_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_2335_),
    .B(_1206_),
    .Y(_2336_));
 sky130_fd_sc_hd__nand2_1 _5712_ (.A(_2336_),
    .B(_1102_),
    .Y(_2337_));
 sky130_fd_sc_hd__nand2_1 _5713_ (.A(_2337_),
    .B(_2316_),
    .Y(_2338_));
 sky130_fd_sc_hd__a21oi_1 _5714_ (.A1(_0787_),
    .A2(\BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2339_));
 sky130_fd_sc_hd__nand2_1 _5715_ (.A(_2338_),
    .B(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__nand2_2 _5716_ (.A(_2340_),
    .B(_2311_),
    .Y(_2341_));
 sky130_fd_sc_hd__o21ai_1 _5717_ (.A1(\BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(\BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_1622_),
    .Y(_2342_));
 sky130_fd_sc_hd__o211a_1 _5718_ (.A1(\BitStream_buffer.BitStream_buffer_output[5] ),
    .A2(_2342_),
    .B1(_1310_),
    .C1(_1414_),
    .X(_2343_));
 sky130_fd_sc_hd__a21o_1 _5719_ (.A1(_2315_),
    .A2(_2325_),
    .B1(_2312_),
    .X(_2344_));
 sky130_fd_sc_hd__o21bai_4 _5720_ (.A1(_2343_),
    .A2(_2318_),
    .B1_N(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__nor2_2 _5721_ (.A(\BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\BitStream_buffer.BitStream_buffer_valid_n ),
    .Y(_2346_));
 sky130_fd_sc_hd__nand3_1 _5722_ (.A(_2341_),
    .B(_2345_),
    .C(_2346_),
    .Y(_2347_));
 sky130_fd_sc_hd__nor2_1 _5723_ (.A(_2329_),
    .B(_2347_),
    .Y(_2348_));
 sky130_fd_sc_hd__inv_2 _5724_ (.A(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__nor2_1 _5725_ (.A(\BitStream_buffer.BitStream_buffer_output[5] ),
    .B(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__inv_4 _5726_ (.A(_2345_),
    .Y(_2351_));
 sky130_fd_sc_hd__nor2_1 _5727_ (.A(_2351_),
    .B(_2329_),
    .Y(_2352_));
 sky130_fd_sc_hd__nand2_2 _5728_ (.A(_2341_),
    .B(_2346_),
    .Y(_2353_));
 sky130_fd_sc_hd__nand2_1 _5729_ (.A(_2352_),
    .B(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__nand2_1 _5730_ (.A(_2351_),
    .B(_2326_),
    .Y(_2355_));
 sky130_fd_sc_hd__inv_2 _5731_ (.A(_2355_),
    .Y(_2356_));
 sky130_fd_sc_hd__nand3_1 _5732_ (.A(_2356_),
    .B(_2353_),
    .C(_0894_),
    .Y(_2357_));
 sky130_fd_sc_hd__o21ai_1 _5733_ (.A1(\BitStream_buffer.BitStream_buffer_output[7] ),
    .A2(_2354_),
    .B1(_2357_),
    .Y(_2358_));
 sky130_fd_sc_hd__nor2_1 _5734_ (.A(_2350_),
    .B(_2358_),
    .Y(_2359_));
 sky130_fd_sc_hd__nand3_4 _5735_ (.A(_2341_),
    .B(_2351_),
    .C(_2346_),
    .Y(_2360_));
 sky130_fd_sc_hd__inv_4 _5736_ (.A(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__and3_1 _5737_ (.A(_2361_),
    .B(_1102_),
    .C(_2326_),
    .X(_2362_));
 sky130_fd_sc_hd__inv_2 _5738_ (.A(_2347_),
    .Y(_2363_));
 sky130_fd_sc_hd__and3_1 _5739_ (.A(_2363_),
    .B(_0671_),
    .C(_2326_),
    .X(_2364_));
 sky130_fd_sc_hd__nor2_1 _5740_ (.A(_2362_),
    .B(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(_2361_),
    .B(_2328_),
    .Y(_2366_));
 sky130_fd_sc_hd__nand2_1 _5742_ (.A(_2366_),
    .B(_1726_),
    .Y(_2367_));
 sky130_fd_sc_hd__nor2_1 _5743_ (.A(_2329_),
    .B(_2360_),
    .Y(_2368_));
 sky130_fd_sc_hd__nand2_1 _5744_ (.A(_2368_),
    .B(_1934_),
    .Y(_2369_));
 sky130_fd_sc_hd__nand2_1 _5745_ (.A(_2367_),
    .B(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__nor2_2 _5746_ (.A(_2345_),
    .B(_2329_),
    .Y(_2371_));
 sky130_fd_sc_hd__nand2_1 _5747_ (.A(_2370_),
    .B(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__nand3_2 _5748_ (.A(_2359_),
    .B(_2365_),
    .C(_2372_),
    .Y(_2373_));
 sky130_fd_sc_hd__nand2_2 _5749_ (.A(_2373_),
    .B(_2607_),
    .Y(_2374_));
 sky130_fd_sc_hd__inv_2 _5750_ (.A(_2374_),
    .Y(_2375_));
 sky130_fd_sc_hd__or2_1 _5751_ (.A(_2310_),
    .B(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__a311o_1 _5752_ (.A1(_2353_),
    .A2(_2327_),
    .A3(_2345_),
    .B1(_2608_),
    .C1(_2319_),
    .X(_2377_));
 sky130_fd_sc_hd__nand2_1 _5753_ (.A(_2377_),
    .B(_2310_),
    .Y(_2378_));
 sky130_fd_sc_hd__nor2_1 _5754_ (.A(net18),
    .B(_2606_),
    .Y(_2379_));
 sky130_fd_sc_hd__nand2_1 _5755_ (.A(_2366_),
    .B(\BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2380_));
 sky130_fd_sc_hd__buf_6 _5756_ (.A(_2368_),
    .X(_2381_));
 sky130_fd_sc_hd__nand2_1 _5757_ (.A(_2381_),
    .B(\BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2382_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(_2380_),
    .B(_2382_),
    .Y(_2383_));
 sky130_fd_sc_hd__nand2_1 _5759_ (.A(_2370_),
    .B(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__o21ai_1 _5760_ (.A1(_2329_),
    .A2(_2360_),
    .B1(\BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2385_));
 sky130_fd_sc_hd__nand2_1 _5761_ (.A(_2381_),
    .B(\BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2386_));
 sky130_fd_sc_hd__nand2_1 _5762_ (.A(_2385_),
    .B(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__o21ai_1 _5763_ (.A1(_2329_),
    .A2(_2360_),
    .B1(_1622_),
    .Y(_2388_));
 sky130_fd_sc_hd__nand3_1 _5764_ (.A(_2361_),
    .B(_1830_),
    .C(_2328_),
    .Y(_2389_));
 sky130_fd_sc_hd__nand2_1 _5765_ (.A(_2388_),
    .B(_2389_),
    .Y(_2390_));
 sky130_fd_sc_hd__nand2_1 _5766_ (.A(_2387_),
    .B(_2390_),
    .Y(_2391_));
 sky130_fd_sc_hd__nand3_1 _5767_ (.A(_2384_),
    .B(_2391_),
    .C(_2371_),
    .Y(_2392_));
 sky130_fd_sc_hd__and2_1 _5768_ (.A(_2361_),
    .B(_2326_),
    .X(_2393_));
 sky130_fd_sc_hd__nor2_1 _5769_ (.A(\BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2394_));
 sky130_fd_sc_hd__inv_2 _5770_ (.A(_2394_),
    .Y(_2395_));
 sky130_fd_sc_hd__nand2_1 _5771_ (.A(\BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2396_));
 sky130_fd_sc_hd__nand2_1 _5772_ (.A(_2395_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__nand2_1 _5773_ (.A(_2393_),
    .B(_2397_),
    .Y(_2398_));
 sky130_fd_sc_hd__xnor2_1 _5774_ (.A(\BitStream_buffer.BitStream_buffer_output[14] ),
    .B(\BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2399_));
 sky130_fd_sc_hd__nand3_1 _5775_ (.A(_2363_),
    .B(_2326_),
    .C(_2399_),
    .Y(_2400_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(_2398_),
    .B(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__xor2_1 _5777_ (.A(\BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\BitStream_buffer.BitStream_buffer_output[11] ),
    .X(_2402_));
 sky130_fd_sc_hd__nand2_1 _5778_ (.A(_2356_),
    .B(_2353_),
    .Y(_2403_));
 sky130_fd_sc_hd__nor2_2 _5779_ (.A(\BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2404_));
 sky130_fd_sc_hd__inv_2 _5780_ (.A(_2404_),
    .Y(_2405_));
 sky130_fd_sc_hd__nand2_1 _5781_ (.A(\BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2406_));
 sky130_fd_sc_hd__nand2_1 _5782_ (.A(_2405_),
    .B(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__nand3_1 _5783_ (.A(_2352_),
    .B(_2353_),
    .C(_2407_),
    .Y(_2408_));
 sky130_fd_sc_hd__nand2_1 _5784_ (.A(\BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2409_));
 sky130_fd_sc_hd__nand2_1 _5785_ (.A(_2321_),
    .B(_2409_),
    .Y(_2410_));
 sky130_fd_sc_hd__nand2_1 _5786_ (.A(_2348_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__o211ai_1 _5787_ (.A1(_2402_),
    .A2(_2403_),
    .B1(_2408_),
    .C1(_2411_),
    .Y(_2412_));
 sky130_fd_sc_hd__nor2_1 _5788_ (.A(_2401_),
    .B(_2412_),
    .Y(_2413_));
 sky130_fd_sc_hd__nand2_1 _5789_ (.A(_2392_),
    .B(_2413_),
    .Y(_2414_));
 sky130_fd_sc_hd__buf_4 _5790_ (.A(_2607_),
    .X(_2415_));
 sky130_fd_sc_hd__nand3_1 _5791_ (.A(_2414_),
    .B(_2415_),
    .C(_2373_),
    .Y(_2416_));
 sky130_fd_sc_hd__nor2_2 _5792_ (.A(net17),
    .B(_2605_),
    .Y(_2417_));
 sky130_fd_sc_hd__a22o_1 _5793_ (.A1(_2375_),
    .A2(_2379_),
    .B1(_2416_),
    .B2(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__nand2_1 _5794_ (.A(_2414_),
    .B(_2607_),
    .Y(_2419_));
 sky130_fd_sc_hd__nand2_1 _5795_ (.A(_2419_),
    .B(_2374_),
    .Y(_2420_));
 sky130_fd_sc_hd__a32o_1 _5796_ (.A1(_2307_),
    .A2(_2376_),
    .A3(_2378_),
    .B1(_2418_),
    .B2(_2420_),
    .X(net20));
 sky130_fd_sc_hd__a31o_1 _5797_ (.A1(_2308_),
    .A2(net18),
    .A3(_2309_),
    .B1(_2606_),
    .X(_2421_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_2370_),
    .B(_2390_),
    .Y(_2422_));
 sky130_fd_sc_hd__o21ai_1 _5799_ (.A1(_2329_),
    .A2(_2360_),
    .B1(_1518_),
    .Y(_2423_));
 sky130_fd_sc_hd__nand3_1 _5800_ (.A(_2361_),
    .B(_1726_),
    .C(_2328_),
    .Y(_2424_));
 sky130_fd_sc_hd__nand2_1 _5801_ (.A(_2423_),
    .B(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__nand2_1 _5802_ (.A(_2422_),
    .B(_2425_),
    .Y(_2426_));
 sky130_fd_sc_hd__o21ai_1 _5803_ (.A1(_2329_),
    .A2(_2360_),
    .B1(\BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2427_));
 sky130_fd_sc_hd__nand2_1 _5804_ (.A(_2381_),
    .B(\BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2428_));
 sky130_fd_sc_hd__nand2_1 _5805_ (.A(_2427_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__nand3_1 _5806_ (.A(_2370_),
    .B(_2429_),
    .C(_2390_),
    .Y(_2430_));
 sky130_fd_sc_hd__nand3_1 _5807_ (.A(_2426_),
    .B(_2430_),
    .C(_2371_),
    .Y(_2431_));
 sky130_fd_sc_hd__nor2_1 _5808_ (.A(\BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2395_),
    .Y(_2432_));
 sky130_fd_sc_hd__nor2_1 _5809_ (.A(_0894_),
    .B(_2394_),
    .Y(_2433_));
 sky130_fd_sc_hd__o21ai_1 _5810_ (.A1(_2432_),
    .A2(_2433_),
    .B1(_2393_),
    .Y(_2434_));
 sky130_fd_sc_hd__nor2_1 _5811_ (.A(_1310_),
    .B(_2320_),
    .Y(_2435_));
 sky130_fd_sc_hd__o21ai_1 _5812_ (.A1(_2322_),
    .A2(_2435_),
    .B1(_2348_),
    .Y(_2436_));
 sky130_fd_sc_hd__nand2_1 _5813_ (.A(_2434_),
    .B(_2436_),
    .Y(_2437_));
 sky130_fd_sc_hd__and2_1 _5814_ (.A(_2313_),
    .B(\BitStream_buffer.BitStream_buffer_output[13] ),
    .X(_2438_));
 sky130_fd_sc_hd__nor2_1 _5815_ (.A(_2314_),
    .B(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__nor2_1 _5816_ (.A(_1102_),
    .B(_2404_),
    .Y(_2440_));
 sky130_fd_sc_hd__nor2_1 _5817_ (.A(\BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2405_),
    .Y(_2441_));
 sky130_fd_sc_hd__inv_2 _5818_ (.A(_2354_),
    .Y(_2442_));
 sky130_fd_sc_hd__o21ai_1 _5819_ (.A1(_2440_),
    .A2(_2441_),
    .B1(_2442_),
    .Y(_2443_));
 sky130_fd_sc_hd__o21ai_1 _5820_ (.A1(_2403_),
    .A2(_2439_),
    .B1(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__nor2_1 _5821_ (.A(_2437_),
    .B(_2444_),
    .Y(_2445_));
 sky130_fd_sc_hd__nand2_1 _5822_ (.A(_2431_),
    .B(_2445_),
    .Y(_2446_));
 sky130_fd_sc_hd__nand2_1 _5823_ (.A(_2446_),
    .B(_2415_),
    .Y(_2447_));
 sky130_fd_sc_hd__nand2_2 _5824_ (.A(_2447_),
    .B(_2419_),
    .Y(_2448_));
 sky130_fd_sc_hd__nand3_1 _5825_ (.A(_2446_),
    .B(_2415_),
    .C(_2414_),
    .Y(_2449_));
 sky130_fd_sc_hd__nand3_1 _5826_ (.A(_2448_),
    .B(_2417_),
    .C(_2449_),
    .Y(_2450_));
 sky130_fd_sc_hd__o21ai_2 _5827_ (.A1(_2419_),
    .A2(_2421_),
    .B1(_2450_),
    .Y(net21));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_2449_),
    .B(_2375_),
    .Y(_2451_));
 sky130_fd_sc_hd__nand2_1 _5829_ (.A(_2451_),
    .B(_2448_),
    .Y(_2452_));
 sky130_fd_sc_hd__nor2_1 _5830_ (.A(_2387_),
    .B(_2383_),
    .Y(_2453_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(_2381_),
    .B(\BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2454_));
 sky130_fd_sc_hd__o21ai_1 _5832_ (.A1(_1414_),
    .A2(_2381_),
    .B1(_2454_),
    .Y(_2455_));
 sky130_fd_sc_hd__nand3_1 _5833_ (.A(_2453_),
    .B(_2425_),
    .C(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hd__nand3_1 _5834_ (.A(_2370_),
    .B(_2390_),
    .C(_2425_),
    .Y(_2457_));
 sky130_fd_sc_hd__nand2_1 _5835_ (.A(_2368_),
    .B(_1622_),
    .Y(_2458_));
 sky130_fd_sc_hd__o21ai_1 _5836_ (.A1(\BitStream_buffer.BitStream_buffer_output[6] ),
    .A2(_2381_),
    .B1(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_2457_),
    .B(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__nand3_1 _5838_ (.A(_2456_),
    .B(_2460_),
    .C(_2371_),
    .Y(_2461_));
 sky130_fd_sc_hd__or2_1 _5839_ (.A(\BitStream_buffer.BitStream_buffer_output[12] ),
    .B(_2432_),
    .X(_2462_));
 sky130_fd_sc_hd__nand2_1 _5840_ (.A(_2432_),
    .B(\BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2463_));
 sky130_fd_sc_hd__and3_1 _5841_ (.A(_2393_),
    .B(_2462_),
    .C(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__or2_1 _5842_ (.A(_1206_),
    .B(_2322_),
    .X(_2465_));
 sky130_fd_sc_hd__nor2_1 _5843_ (.A(_2321_),
    .B(_2405_),
    .Y(_2466_));
 sky130_fd_sc_hd__inv_2 _5844_ (.A(_2466_),
    .Y(_2467_));
 sky130_fd_sc_hd__nand2_1 _5845_ (.A(_2465_),
    .B(_2467_),
    .Y(_2468_));
 sky130_fd_sc_hd__mux2_1 _5846_ (.A0(\BitStream_buffer.BitStream_buffer_output[10] ),
    .A1(_2397_),
    .S(_2404_),
    .X(_2469_));
 sky130_fd_sc_hd__a22o_1 _5847_ (.A1(_2348_),
    .A2(_2468_),
    .B1(_2442_),
    .B2(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__nor2_1 _5848_ (.A(_2464_),
    .B(_2470_),
    .Y(_2471_));
 sky130_fd_sc_hd__a21oi_2 _5849_ (.A1(_2461_),
    .A2(_2471_),
    .B1(_2608_),
    .Y(_2472_));
 sky130_fd_sc_hd__nand2_1 _5850_ (.A(_2452_),
    .B(_2472_),
    .Y(_2473_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_2461_),
    .B(_2471_),
    .Y(_2474_));
 sky130_fd_sc_hd__nand2_1 _5852_ (.A(_2474_),
    .B(_2415_),
    .Y(_2475_));
 sky130_fd_sc_hd__nand3_1 _5853_ (.A(_2451_),
    .B(_2448_),
    .C(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__nand2_1 _5854_ (.A(_2473_),
    .B(_2476_),
    .Y(_2477_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_2477_),
    .B(_2417_),
    .Y(_2478_));
 sky130_fd_sc_hd__or2_1 _5856_ (.A(_2421_),
    .B(_2447_),
    .X(_2479_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(_2478_),
    .B(_2479_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_1 _5858_ (.A(net20),
    .B(net21),
    .Y(_2480_));
 sky130_fd_sc_hd__inv_2 _5859_ (.A(_2480_),
    .Y(_2481_));
 sky130_fd_sc_hd__nand2_1 _5860_ (.A(net22),
    .B(_2481_),
    .Y(_2482_));
 sky130_fd_sc_hd__nand3_1 _5861_ (.A(_2478_),
    .B(_2480_),
    .C(_2479_),
    .Y(_2483_));
 sky130_fd_sc_hd__nand3_1 _5862_ (.A(_2482_),
    .B(_2307_),
    .C(_2483_),
    .Y(_2484_));
 sky130_fd_sc_hd__inv_2 _5863_ (.A(_2484_),
    .Y(\exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__or3_1 _5864_ (.A(_2608_),
    .B(_2310_),
    .C(_2353_),
    .X(_2485_));
 sky130_fd_sc_hd__inv_2 _5865_ (.A(_2485_),
    .Y(\BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__or3_1 _5866_ (.A(_2608_),
    .B(_2310_),
    .C(_2345_),
    .X(_2486_));
 sky130_fd_sc_hd__inv_2 _5867_ (.A(_2486_),
    .Y(\BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__or3_1 _5868_ (.A(_2608_),
    .B(_2310_),
    .C(_2327_),
    .X(_2487_));
 sky130_fd_sc_hd__inv_2 _5869_ (.A(_2487_),
    .Y(\BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__nand2_1 _5870_ (.A(_2459_),
    .B(_2425_),
    .Y(_2488_));
 sky130_fd_sc_hd__nor2_1 _5871_ (.A(_2422_),
    .B(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__nand2_1 _5872_ (.A(_2381_),
    .B(\BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2490_));
 sky130_fd_sc_hd__o21ai_2 _5873_ (.A1(_1310_),
    .A2(_2381_),
    .B1(_2490_),
    .Y(_2491_));
 sky130_fd_sc_hd__nand2_1 _5874_ (.A(_2489_),
    .B(_2491_),
    .Y(_2492_));
 sky130_fd_sc_hd__nor2_1 _5875_ (.A(_2429_),
    .B(_2455_),
    .Y(_2493_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_2493_),
    .B(_2453_),
    .Y(_2494_));
 sky130_fd_sc_hd__inv_2 _5877_ (.A(_2491_),
    .Y(_2495_));
 sky130_fd_sc_hd__nand2_1 _5878_ (.A(_2494_),
    .B(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__nand3_1 _5879_ (.A(_2492_),
    .B(_2496_),
    .C(_2371_),
    .Y(_2497_));
 sky130_fd_sc_hd__nor2_1 _5880_ (.A(_1102_),
    .B(_2467_),
    .Y(_2498_));
 sky130_fd_sc_hd__nor2_1 _5881_ (.A(\BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2466_),
    .Y(_2499_));
 sky130_fd_sc_hd__nand2_1 _5882_ (.A(_2404_),
    .B(_2394_),
    .Y(_2500_));
 sky130_fd_sc_hd__xor2_1 _5883_ (.A(\BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__o32a_1 _5884_ (.A1(_2498_),
    .A2(_2499_),
    .A3(_2349_),
    .B1(_2354_),
    .B2(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__nand2_1 _5885_ (.A(_2497_),
    .B(_2502_),
    .Y(_2503_));
 sky130_fd_sc_hd__nand2_2 _5886_ (.A(_2503_),
    .B(_2415_),
    .Y(_2504_));
 sky130_fd_sc_hd__nor2_1 _5887_ (.A(_2448_),
    .B(_2472_),
    .Y(_2505_));
 sky130_fd_sc_hd__nor2_1 _5888_ (.A(_2504_),
    .B(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__nand2_1 _5889_ (.A(_2504_),
    .B(_2475_),
    .Y(_2507_));
 sky130_fd_sc_hd__nor2_1 _5890_ (.A(_2448_),
    .B(_2507_),
    .Y(_2508_));
 sky130_fd_sc_hd__o21a_1 _5891_ (.A1(_2506_),
    .A2(_2508_),
    .B1(_2374_),
    .X(_2509_));
 sky130_fd_sc_hd__nor2_1 _5892_ (.A(_2416_),
    .B(_2447_),
    .Y(_2510_));
 sky130_fd_sc_hd__nand2_1 _5893_ (.A(_2472_),
    .B(_2510_),
    .Y(_2511_));
 sky130_fd_sc_hd__nor2_1 _5894_ (.A(_2504_),
    .B(_2511_),
    .Y(_2512_));
 sky130_fd_sc_hd__and2_1 _5895_ (.A(_2511_),
    .B(_2504_),
    .X(_2513_));
 sky130_fd_sc_hd__o21ai_1 _5896_ (.A1(_2512_),
    .A2(_2513_),
    .B1(_2375_),
    .Y(_2514_));
 sky130_fd_sc_hd__nand2_1 _5897_ (.A(_2514_),
    .B(_2417_),
    .Y(_2515_));
 sky130_fd_sc_hd__inv_2 _5898_ (.A(_2421_),
    .Y(_2516_));
 sky130_fd_sc_hd__nand2_1 _5899_ (.A(_2474_),
    .B(_2516_),
    .Y(_2517_));
 sky130_fd_sc_hd__o21ai_2 _5900_ (.A1(_2509_),
    .A2(_2515_),
    .B1(_2517_),
    .Y(net23));
 sky130_fd_sc_hd__nand2_1 _5901_ (.A(_2508_),
    .B(_2374_),
    .Y(_2518_));
 sky130_fd_sc_hd__o21ai_1 _5902_ (.A1(_2504_),
    .A2(_2511_),
    .B1(_2375_),
    .Y(_2519_));
 sky130_fd_sc_hd__nand2_1 _5903_ (.A(_2518_),
    .B(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__nand3_1 _5904_ (.A(_2493_),
    .B(_2453_),
    .C(_2495_),
    .Y(_2521_));
 sky130_fd_sc_hd__a21oi_2 _5905_ (.A1(_2381_),
    .A2(_1414_),
    .B1(_1206_),
    .Y(_2522_));
 sky130_fd_sc_hd__inv_2 _5906_ (.A(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(_2521_),
    .B(_2523_),
    .Y(_2524_));
 sky130_fd_sc_hd__nand3_1 _5908_ (.A(_2489_),
    .B(_2495_),
    .C(_2522_),
    .Y(_2525_));
 sky130_fd_sc_hd__nand3_1 _5909_ (.A(_2524_),
    .B(_2525_),
    .C(_2371_),
    .Y(_2526_));
 sky130_fd_sc_hd__nor2_1 _5910_ (.A(_2397_),
    .B(_2467_),
    .Y(_2527_));
 sky130_fd_sc_hd__a211o_1 _5911_ (.A1(_0998_),
    .A2(_2467_),
    .B1(_2527_),
    .C1(_2349_),
    .X(_2528_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(_2526_),
    .B(_2528_),
    .Y(_2529_));
 sky130_fd_sc_hd__nand2_1 _5913_ (.A(_2529_),
    .B(_2415_),
    .Y(_2530_));
 sky130_fd_sc_hd__nand2_1 _5914_ (.A(_2520_),
    .B(_2530_),
    .Y(_2531_));
 sky130_fd_sc_hd__inv_2 _5915_ (.A(_2530_),
    .Y(_2532_));
 sky130_fd_sc_hd__nand3_1 _5916_ (.A(_2518_),
    .B(_2519_),
    .C(_2532_),
    .Y(_2533_));
 sky130_fd_sc_hd__nand3_1 _5917_ (.A(_2531_),
    .B(_2533_),
    .C(_2417_),
    .Y(_2534_));
 sky130_fd_sc_hd__nand2_1 _5918_ (.A(_2503_),
    .B(_2516_),
    .Y(_2535_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_2534_),
    .B(_2535_),
    .Y(net24));
 sky130_fd_sc_hd__nand3_1 _5920_ (.A(_2529_),
    .B(_2415_),
    .C(_2503_),
    .Y(_2536_));
 sky130_fd_sc_hd__inv_2 _5921_ (.A(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__nor3_1 _5922_ (.A(_2447_),
    .B(_2416_),
    .C(_2475_),
    .Y(_2538_));
 sky130_fd_sc_hd__nand2_1 _5923_ (.A(_2537_),
    .B(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(_2328_),
    .B(_2351_),
    .Y(_2540_));
 sky130_fd_sc_hd__nor2_1 _5925_ (.A(_2522_),
    .B(_2491_),
    .Y(_2541_));
 sky130_fd_sc_hd__nand2_1 _5926_ (.A(_2489_),
    .B(_2541_),
    .Y(_2542_));
 sky130_fd_sc_hd__o21ai_2 _5927_ (.A1(_1310_),
    .A2(_2366_),
    .B1(_1102_),
    .Y(_2543_));
 sky130_fd_sc_hd__inv_2 _5928_ (.A(_2543_),
    .Y(_2544_));
 sky130_fd_sc_hd__nand2_1 _5929_ (.A(_2542_),
    .B(_2544_),
    .Y(_2545_));
 sky130_fd_sc_hd__nand3_1 _5930_ (.A(_2489_),
    .B(_2541_),
    .C(_2543_),
    .Y(_2546_));
 sky130_fd_sc_hd__nand2_1 _5931_ (.A(_2545_),
    .B(_2546_),
    .Y(_2547_));
 sky130_fd_sc_hd__nor2_1 _5932_ (.A(_2540_),
    .B(_2547_),
    .Y(_2548_));
 sky130_fd_sc_hd__nand2_1 _5933_ (.A(_2548_),
    .B(_2415_),
    .Y(_2549_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(_2539_),
    .B(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__inv_2 _5935_ (.A(_2549_),
    .Y(_2551_));
 sky130_fd_sc_hd__nand3_1 _5936_ (.A(_2537_),
    .B(_2538_),
    .C(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(_2550_),
    .B(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__nand2_1 _5938_ (.A(_2553_),
    .B(_2375_),
    .Y(_2554_));
 sky130_fd_sc_hd__nand3_1 _5939_ (.A(_2505_),
    .B(_2530_),
    .C(_2504_),
    .Y(_2555_));
 sky130_fd_sc_hd__nand2b_1 _5940_ (.A_N(_2547_),
    .B(_2371_),
    .Y(_2556_));
 sky130_fd_sc_hd__nor2_1 _5941_ (.A(_2608_),
    .B(_2556_),
    .Y(_2557_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_2555_),
    .B(_2557_),
    .Y(_2558_));
 sky130_fd_sc_hd__o21ai_1 _5943_ (.A1(_2548_),
    .A2(_2529_),
    .B1(_2415_),
    .Y(_2559_));
 sky130_fd_sc_hd__nand2_1 _5944_ (.A(_2508_),
    .B(_2559_),
    .Y(_2560_));
 sky130_fd_sc_hd__nand2_1 _5945_ (.A(_2558_),
    .B(_2560_),
    .Y(_2561_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(_2561_),
    .B(_2374_),
    .Y(_2562_));
 sky130_fd_sc_hd__nand3_1 _5947_ (.A(_2554_),
    .B(_2417_),
    .C(_2562_),
    .Y(_2563_));
 sky130_fd_sc_hd__nand2_1 _5948_ (.A(_2529_),
    .B(_2516_),
    .Y(_2564_));
 sky130_fd_sc_hd__nand2_1 _5949_ (.A(_2563_),
    .B(_2564_),
    .Y(net25));
 sky130_fd_sc_hd__nand3_1 _5950_ (.A(_2512_),
    .B(_2532_),
    .C(_2557_),
    .Y(_2565_));
 sky130_fd_sc_hd__or2_1 _5951_ (.A(_2543_),
    .B(_2542_),
    .X(_2566_));
 sky130_fd_sc_hd__nand2_1 _5952_ (.A(_2566_),
    .B(_2381_),
    .Y(_2567_));
 sky130_fd_sc_hd__inv_2 _5953_ (.A(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__nand2_1 _5954_ (.A(_2568_),
    .B(_2415_),
    .Y(_2569_));
 sky130_fd_sc_hd__nand2_1 _5955_ (.A(_2565_),
    .B(_2569_),
    .Y(_2570_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_2570_),
    .B(_2375_),
    .Y(_2571_));
 sky130_fd_sc_hd__inv_2 _5957_ (.A(_2569_),
    .Y(_2572_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_2560_),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__nor2_1 _5959_ (.A(_2377_),
    .B(_2373_),
    .Y(_2574_));
 sky130_fd_sc_hd__nand2_1 _5960_ (.A(_2573_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__nand2_1 _5961_ (.A(_2571_),
    .B(_2575_),
    .Y(_2576_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(_2576_),
    .B(_2417_),
    .Y(_2577_));
 sky130_fd_sc_hd__a211o_1 _5963_ (.A1(net18),
    .A2(_2310_),
    .B1(_2606_),
    .C1(_2556_),
    .X(_2578_));
 sky130_fd_sc_hd__nand2_1 _5964_ (.A(_2577_),
    .B(_2578_),
    .Y(net26));
 sky130_fd_sc_hd__a211o_1 _5965_ (.A1(net18),
    .A2(_2310_),
    .B1(_2606_),
    .C1(_2567_),
    .X(_2579_));
 sky130_fd_sc_hd__a21bo_1 _5966_ (.A1(_2417_),
    .A2(_2574_),
    .B1_N(_2579_),
    .X(net27));
 sky130_fd_sc_hd__buf_1 _5967_ (.A(clk),
    .X(_2580_));
 sky130_fd_sc_hd__buf_1 _5968_ (.A(clknet_1_0__leaf__2580_),
    .X(_2581_));
 sky130_fd_sc_hd__buf_1 _5969_ (.A(clknet_1_0__leaf__2581_),
    .X(_2582_));
 sky130_fd_sc_hd__inv_2 _5970__72 (.A(clknet_1_1__leaf__2582_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _5971__73 (.A(clknet_1_1__leaf__2582_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _5972__74 (.A(clknet_1_1__leaf__2582_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _5973__75 (.A(clknet_1_0__leaf__2582_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _5974__76 (.A(clknet_1_1__leaf__2582_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _5975__77 (.A(clknet_1_0__leaf__2582_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _5976__78 (.A(clknet_1_0__leaf__2582_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _5977__79 (.A(clknet_1_0__leaf__2582_),
    .Y(net115));
 sky130_fd_sc_hd__inv_2 _5978__80 (.A(clknet_1_0__leaf__2582_),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _5979__81 (.A(clknet_1_0__leaf__2582_),
    .Y(net117));
 sky130_fd_sc_hd__buf_1 _5980_ (.A(clknet_1_0__leaf__2581_),
    .X(_2583_));
 sky130_fd_sc_hd__inv_2 _5981__82 (.A(clknet_1_0__leaf__2583_),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _5982__83 (.A(clknet_1_1__leaf__2583_),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _5983__84 (.A(clknet_1_0__leaf__2583_),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _5984__85 (.A(clknet_1_0__leaf__2583_),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _5985__86 (.A(clknet_1_0__leaf__2583_),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _5986__87 (.A(clknet_1_1__leaf__2583_),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _5987__88 (.A(clknet_1_1__leaf__2583_),
    .Y(net124));
 sky130_fd_sc_hd__inv_2 _5988__89 (.A(clknet_1_1__leaf__2583_),
    .Y(net125));
 sky130_fd_sc_hd__inv_2 _5989__90 (.A(clknet_1_1__leaf__2583_),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _5990__91 (.A(clknet_1_1__leaf__2583_),
    .Y(net127));
 sky130_fd_sc_hd__buf_1 _5991_ (.A(clknet_1_0__leaf__2581_),
    .X(_2584_));
 sky130_fd_sc_hd__inv_2 _5992__92 (.A(clknet_1_0__leaf__2584_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _5993__93 (.A(clknet_1_0__leaf__2584_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _5994__94 (.A(clknet_1_0__leaf__2584_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _5995__95 (.A(clknet_1_0__leaf__2584_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _5996__96 (.A(clknet_1_1__leaf__2584_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _5997__97 (.A(clknet_1_1__leaf__2584_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _5998__98 (.A(clknet_1_1__leaf__2584_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _5999__99 (.A(clknet_1_1__leaf__2584_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _6000__100 (.A(clknet_1_1__leaf__2584_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _6001__101 (.A(clknet_1_1__leaf__2584_),
    .Y(net137));
 sky130_fd_sc_hd__buf_1 _6002_ (.A(clknet_1_0__leaf__2581_),
    .X(_2585_));
 sky130_fd_sc_hd__inv_2 _6003__102 (.A(clknet_1_0__leaf__2585_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _6004__103 (.A(clknet_1_0__leaf__2585_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _6005__104 (.A(clknet_1_0__leaf__2585_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _6006__105 (.A(clknet_1_0__leaf__2585_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _6007__106 (.A(clknet_1_0__leaf__2585_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _6008__107 (.A(clknet_1_0__leaf__2585_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _6009__108 (.A(clknet_1_1__leaf__2585_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _6010__109 (.A(clknet_1_1__leaf__2585_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _6011__110 (.A(clknet_1_1__leaf__2585_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _6012__111 (.A(clknet_1_1__leaf__2585_),
    .Y(net147));
 sky130_fd_sc_hd__buf_1 _6013_ (.A(clknet_1_1__leaf__2581_),
    .X(_2586_));
 sky130_fd_sc_hd__inv_2 _6014__112 (.A(clknet_1_0__leaf__2586_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _6015__113 (.A(clknet_1_0__leaf__2586_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _6016__114 (.A(clknet_1_0__leaf__2586_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _6017__115 (.A(clknet_1_0__leaf__2586_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _6018__116 (.A(clknet_1_1__leaf__2586_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _6019__117 (.A(clknet_1_1__leaf__2586_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _6020__118 (.A(clknet_1_1__leaf__2586_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _6021__119 (.A(clknet_1_1__leaf__2586_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _6022__120 (.A(clknet_1_1__leaf__2586_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _6023__121 (.A(clknet_1_1__leaf__2586_),
    .Y(net157));
 sky130_fd_sc_hd__buf_1 _6024_ (.A(clknet_1_1__leaf__2581_),
    .X(_2587_));
 sky130_fd_sc_hd__inv_2 _6025__122 (.A(clknet_1_1__leaf__2587_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _6026__123 (.A(clknet_1_0__leaf__2587_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _6027__124 (.A(clknet_1_0__leaf__2587_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _6028__125 (.A(clknet_1_0__leaf__2587_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _6029__126 (.A(clknet_1_0__leaf__2587_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _6030__127 (.A(clknet_1_0__leaf__2587_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _6031__128 (.A(clknet_1_0__leaf__2587_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _6032__129 (.A(clknet_1_1__leaf__2587_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _6033__130 (.A(clknet_1_1__leaf__2587_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _6034__131 (.A(clknet_1_1__leaf__2587_),
    .Y(net167));
 sky130_fd_sc_hd__buf_1 _6035_ (.A(clknet_1_1__leaf__2581_),
    .X(_2588_));
 sky130_fd_sc_hd__inv_2 _6036__132 (.A(clknet_1_0__leaf__2588_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _6037__133 (.A(clknet_1_0__leaf__2588_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _6038__134 (.A(clknet_1_0__leaf__2588_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _6039__135 (.A(clknet_1_0__leaf__2588_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _6040__136 (.A(clknet_1_1__leaf__2588_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _6041__137 (.A(clknet_1_1__leaf__2588_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _6042__138 (.A(clknet_1_1__leaf__2588_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _6043__139 (.A(clknet_1_1__leaf__2588_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _6044__140 (.A(clknet_1_1__leaf__2588_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _6045__141 (.A(clknet_1_1__leaf__2588_),
    .Y(net177));
 sky130_fd_sc_hd__buf_1 _6046_ (.A(clknet_1_1__leaf__2581_),
    .X(_2589_));
 sky130_fd_sc_hd__inv_2 _6047__142 (.A(clknet_1_0__leaf__2589_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _6048__143 (.A(clknet_1_0__leaf__2589_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _6049__144 (.A(clknet_1_0__leaf__2589_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _6050__145 (.A(clknet_1_0__leaf__2589_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _6051__146 (.A(clknet_1_0__leaf__2589_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _6052__147 (.A(clknet_1_1__leaf__2589_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _6053__148 (.A(clknet_1_1__leaf__2589_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _6054__149 (.A(clknet_1_1__leaf__2589_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _6055__150 (.A(clknet_1_1__leaf__2589_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _6056__151 (.A(clknet_1_1__leaf__2589_),
    .Y(net187));
 sky130_fd_sc_hd__buf_1 _6057_ (.A(clknet_1_1__leaf__2581_),
    .X(_2590_));
 sky130_fd_sc_hd__inv_2 _6058__152 (.A(clknet_1_1__leaf__2590_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _6059__153 (.A(clknet_1_1__leaf__2590_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _6060__154 (.A(clknet_1_1__leaf__2590_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _6061__155 (.A(clknet_1_0__leaf__2590_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _6062__156 (.A(clknet_1_0__leaf__2590_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _6063__157 (.A(clknet_1_0__leaf__2590_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _6064__158 (.A(clknet_1_0__leaf__2590_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _6065__159 (.A(clknet_1_0__leaf__2590_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _6066__160 (.A(clknet_1_0__leaf__2590_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _6067__161 (.A(clknet_1_1__leaf__2590_),
    .Y(net197));
 sky130_fd_sc_hd__buf_1 _6068_ (.A(clknet_1_1__leaf__2580_),
    .X(_2591_));
 sky130_fd_sc_hd__inv_2 _6069__2 (.A(clknet_1_1__leaf__2591_),
    .Y(net38));
 sky130_fd_sc_hd__inv_2 _6070__3 (.A(clknet_1_1__leaf__2591_),
    .Y(net39));
 sky130_fd_sc_hd__inv_2 _6071__4 (.A(clknet_1_1__leaf__2591_),
    .Y(net40));
 sky130_fd_sc_hd__inv_2 _6072__5 (.A(clknet_1_1__leaf__2591_),
    .Y(net41));
 sky130_fd_sc_hd__inv_2 _6073__6 (.A(clknet_1_1__leaf__2591_),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _6074__7 (.A(clknet_1_0__leaf__2591_),
    .Y(net43));
 sky130_fd_sc_hd__inv_2 _6075__8 (.A(clknet_1_1__leaf__2591_),
    .Y(net44));
 sky130_fd_sc_hd__inv_2 _6076__9 (.A(clknet_1_0__leaf__2591_),
    .Y(net45));
 sky130_fd_sc_hd__inv_2 _6077__10 (.A(clknet_1_0__leaf__2591_),
    .Y(net46));
 sky130_fd_sc_hd__inv_2 _6078__11 (.A(clknet_1_0__leaf__2591_),
    .Y(net47));
 sky130_fd_sc_hd__buf_1 _6079_ (.A(clknet_1_1__leaf__2580_),
    .X(_2592_));
 sky130_fd_sc_hd__inv_2 _6080__12 (.A(clknet_1_0__leaf__2592_),
    .Y(net48));
 sky130_fd_sc_hd__inv_2 _6081__13 (.A(clknet_1_0__leaf__2592_),
    .Y(net49));
 sky130_fd_sc_hd__inv_2 _6082__14 (.A(clknet_1_0__leaf__2592_),
    .Y(net50));
 sky130_fd_sc_hd__inv_2 _6083__15 (.A(clknet_1_0__leaf__2592_),
    .Y(net51));
 sky130_fd_sc_hd__inv_2 _6084__16 (.A(clknet_1_0__leaf__2592_),
    .Y(net52));
 sky130_fd_sc_hd__inv_2 _6085__17 (.A(clknet_1_0__leaf__2592_),
    .Y(net53));
 sky130_fd_sc_hd__inv_2 _6086__18 (.A(clknet_1_1__leaf__2592_),
    .Y(net54));
 sky130_fd_sc_hd__inv_2 _6087__19 (.A(clknet_1_1__leaf__2592_),
    .Y(net55));
 sky130_fd_sc_hd__inv_2 _6088__20 (.A(clknet_1_1__leaf__2592_),
    .Y(net56));
 sky130_fd_sc_hd__inv_2 _6089__21 (.A(clknet_1_1__leaf__2592_),
    .Y(net57));
 sky130_fd_sc_hd__buf_1 _6090_ (.A(clknet_1_1__leaf__2580_),
    .X(_2593_));
 sky130_fd_sc_hd__inv_2 _6091__22 (.A(clknet_1_1__leaf__2593_),
    .Y(net58));
 sky130_fd_sc_hd__inv_2 _6092__23 (.A(clknet_1_1__leaf__2593_),
    .Y(net59));
 sky130_fd_sc_hd__inv_2 _6093__24 (.A(clknet_1_1__leaf__2593_),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 _6094__25 (.A(clknet_1_1__leaf__2593_),
    .Y(net61));
 sky130_fd_sc_hd__inv_2 _6095__26 (.A(clknet_1_0__leaf__2593_),
    .Y(net62));
 sky130_fd_sc_hd__inv_2 _6096__27 (.A(clknet_1_0__leaf__2593_),
    .Y(net63));
 sky130_fd_sc_hd__inv_2 _6097__28 (.A(clknet_1_0__leaf__2593_),
    .Y(net64));
 sky130_fd_sc_hd__inv_2 _6098__29 (.A(clknet_1_0__leaf__2593_),
    .Y(net65));
 sky130_fd_sc_hd__inv_2 _6099__30 (.A(clknet_1_0__leaf__2593_),
    .Y(net66));
 sky130_fd_sc_hd__inv_2 _6100__31 (.A(clknet_1_0__leaf__2593_),
    .Y(net67));
 sky130_fd_sc_hd__buf_1 _6101_ (.A(clknet_1_1__leaf__2580_),
    .X(_2594_));
 sky130_fd_sc_hd__inv_2 _6102__32 (.A(clknet_1_1__leaf__2594_),
    .Y(net68));
 sky130_fd_sc_hd__inv_2 _6103__33 (.A(clknet_1_1__leaf__2594_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _6104__34 (.A(clknet_1_1__leaf__2594_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _6105__35 (.A(clknet_1_1__leaf__2594_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _6106__36 (.A(clknet_1_1__leaf__2594_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _6107__37 (.A(clknet_1_1__leaf__2594_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _6108__38 (.A(clknet_1_0__leaf__2594_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _6109__39 (.A(clknet_1_0__leaf__2594_),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _6110__40 (.A(clknet_1_0__leaf__2594_),
    .Y(net76));
 sky130_fd_sc_hd__inv_2 _6111__41 (.A(clknet_1_0__leaf__2594_),
    .Y(net77));
 sky130_fd_sc_hd__buf_1 _6112_ (.A(clknet_1_0__leaf__2580_),
    .X(_2595_));
 sky130_fd_sc_hd__inv_2 _6113__42 (.A(clknet_1_1__leaf__2595_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _6114__43 (.A(clknet_1_1__leaf__2595_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _6115__44 (.A(clknet_1_1__leaf__2595_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _6116__45 (.A(clknet_1_1__leaf__2595_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _6117__46 (.A(clknet_1_1__leaf__2595_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _6118__47 (.A(clknet_1_0__leaf__2595_),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _6119__48 (.A(clknet_1_0__leaf__2595_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _6120__49 (.A(clknet_1_0__leaf__2595_),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _6121__50 (.A(clknet_1_0__leaf__2595_),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _6122__51 (.A(clknet_1_0__leaf__2595_),
    .Y(net87));
 sky130_fd_sc_hd__buf_1 _6123_ (.A(clknet_1_0__leaf__2580_),
    .X(_2596_));
 sky130_fd_sc_hd__inv_2 _6124__52 (.A(clknet_1_1__leaf__2596_),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _6125__53 (.A(clknet_1_1__leaf__2596_),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _6126__54 (.A(clknet_1_1__leaf__2596_),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _6127__55 (.A(clknet_1_1__leaf__2596_),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _6128__56 (.A(clknet_1_0__leaf__2596_),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _6129__57 (.A(clknet_1_0__leaf__2596_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _6130__58 (.A(clknet_1_0__leaf__2596_),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _6131__59 (.A(clknet_1_0__leaf__2596_),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _6132__60 (.A(clknet_1_0__leaf__2596_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _6133__61 (.A(clknet_1_0__leaf__2596_),
    .Y(net97));
 sky130_fd_sc_hd__buf_1 _6134_ (.A(clknet_1_0__leaf__2580_),
    .X(_2597_));
 sky130_fd_sc_hd__inv_2 _6135__62 (.A(clknet_1_0__leaf__2597_),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _6136__63 (.A(clknet_1_0__leaf__2597_),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _6137__64 (.A(clknet_1_0__leaf__2597_),
    .Y(net100));
 sky130_fd_sc_hd__inv_2 _6138__65 (.A(clknet_1_0__leaf__2597_),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _6139__66 (.A(clknet_1_1__leaf__2597_),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _6140__67 (.A(clknet_1_1__leaf__2597_),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _6141__68 (.A(clknet_1_1__leaf__2597_),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _6142__69 (.A(clknet_1_1__leaf__2597_),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _6143__70 (.A(clknet_1_1__leaf__2597_),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _6144__71 (.A(clknet_1_1__leaf__2597_),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _6145__1 (.A(clknet_1_1__leaf__2581_),
    .Y(net37));
 sky130_fd_sc_hd__dfxtp_1 _6146_ (.CLK(net108),
    .D(_0161_),
    .Q(\BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6147_ (.CLK(net109),
    .D(_0162_),
    .Q(\BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6148_ (.CLK(net110),
    .D(_0163_),
    .Q(\BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6149_ (.CLK(net111),
    .D(_0164_),
    .Q(\BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfxtp_2 _6150_ (.CLK(net112),
    .D(_0165_),
    .Q(\BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfxtp_2 _6151_ (.CLK(net113),
    .D(_0166_),
    .Q(\BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfxtp_2 _6152_ (.CLK(net114),
    .D(_0167_),
    .Q(\BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfxtp_2 _6153_ (.CLK(net115),
    .D(_0168_),
    .Q(\BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfxtp_2 _6154_ (.CLK(net116),
    .D(_0169_),
    .Q(\BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfxtp_2 _6155_ (.CLK(net117),
    .D(_0170_),
    .Q(\BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfxtp_2 _6156_ (.CLK(net118),
    .D(_0171_),
    .Q(\BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfxtp_2 _6157_ (.CLK(net119),
    .D(_0172_),
    .Q(\BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfxtp_2 _6158_ (.CLK(net120),
    .D(_0173_),
    .Q(\BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfxtp_2 _6159_ (.CLK(net121),
    .D(_0174_),
    .Q(\BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfxtp_2 _6160_ (.CLK(net122),
    .D(_0175_),
    .Q(\BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfxtp_2 _6161_ (.CLK(net123),
    .D(_0176_),
    .Q(\BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfxtp_2 _6162_ (.CLK(net124),
    .D(_0177_),
    .Q(\BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfxtp_2 _6163_ (.CLK(net125),
    .D(_0178_),
    .Q(\BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfxtp_2 _6164_ (.CLK(net126),
    .D(_0179_),
    .Q(\BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfxtp_2 _6165_ (.CLK(net127),
    .D(_0180_),
    .Q(\BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfxtp_1 _6166_ (.CLK(net128),
    .D(_0181_),
    .Q(\BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfxtp_1 _6167_ (.CLK(net129),
    .D(_0182_),
    .Q(\BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfxtp_1 _6168_ (.CLK(net130),
    .D(_0183_),
    .Q(\BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfxtp_1 _6169_ (.CLK(net131),
    .D(_0184_),
    .Q(\BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfxtp_1 _6170_ (.CLK(net132),
    .D(_0185_),
    .Q(\BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfxtp_2 _6171_ (.CLK(net133),
    .D(_0186_),
    .Q(\BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfxtp_1 _6172_ (.CLK(net134),
    .D(_0187_),
    .Q(\BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfxtp_2 _6173_ (.CLK(net135),
    .D(_0188_),
    .Q(\BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfxtp_1 _6174_ (.CLK(net136),
    .D(_0189_),
    .Q(\BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfxtp_2 _6175_ (.CLK(net137),
    .D(_0190_),
    .Q(\BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfxtp_1 _6176_ (.CLK(net138),
    .D(_0191_),
    .Q(\BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfxtp_2 _6177_ (.CLK(net139),
    .D(_0192_),
    .Q(\BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfxtp_1 _6178_ (.CLK(net140),
    .D(_0193_),
    .Q(\BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfxtp_2 _6179_ (.CLK(net141),
    .D(_0194_),
    .Q(\BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfxtp_1 _6180_ (.CLK(net142),
    .D(_0195_),
    .Q(\BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfxtp_2 _6181_ (.CLK(net143),
    .D(_0196_),
    .Q(\BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfxtp_2 _6182_ (.CLK(net144),
    .D(_0197_),
    .Q(\BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfxtp_2 _6183_ (.CLK(net145),
    .D(_0198_),
    .Q(\BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfxtp_1 _6184_ (.CLK(net146),
    .D(_0199_),
    .Q(\BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfxtp_1 _6185_ (.CLK(net147),
    .D(_0200_),
    .Q(\BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfxtp_1 _6186_ (.CLK(net148),
    .D(_0201_),
    .Q(\BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfxtp_1 _6187_ (.CLK(net149),
    .D(_0202_),
    .Q(\BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfxtp_1 _6188_ (.CLK(net150),
    .D(_0203_),
    .Q(\BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfxtp_1 _6189_ (.CLK(net151),
    .D(_0204_),
    .Q(\BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfxtp_1 _6190_ (.CLK(net152),
    .D(_0205_),
    .Q(\BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfxtp_1 _6191_ (.CLK(net153),
    .D(_0206_),
    .Q(\BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfxtp_1 _6192_ (.CLK(net154),
    .D(_0207_),
    .Q(\BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfxtp_2 _6193_ (.CLK(net155),
    .D(_0208_),
    .Q(\BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfxtp_2 _6194_ (.CLK(net156),
    .D(_0209_),
    .Q(\BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfxtp_2 _6195_ (.CLK(net157),
    .D(_0210_),
    .Q(\BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfxtp_2 _6196_ (.CLK(net158),
    .D(_0211_),
    .Q(\BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_2 _6197_ (.CLK(net159),
    .D(_0212_),
    .Q(\BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfxtp_2 _6198_ (.CLK(net160),
    .D(_0213_),
    .Q(\BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfxtp_2 _6199_ (.CLK(net161),
    .D(_0214_),
    .Q(\BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfxtp_2 _6200_ (.CLK(net162),
    .D(_0215_),
    .Q(\BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfxtp_2 _6201_ (.CLK(net163),
    .D(_0216_),
    .Q(\BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfxtp_2 _6202_ (.CLK(net164),
    .D(_0217_),
    .Q(\BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfxtp_2 _6203_ (.CLK(net165),
    .D(_0218_),
    .Q(\BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_2 _6204_ (.CLK(net166),
    .D(_0219_),
    .Q(\BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_2 _6205_ (.CLK(net167),
    .D(_0220_),
    .Q(\BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_2 _6206_ (.CLK(net168),
    .D(_0221_),
    .Q(\BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_2 _6207_ (.CLK(net169),
    .D(_0222_),
    .Q(\BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_2 _6208_ (.CLK(net170),
    .D(_0223_),
    .Q(\BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_2 _6209_ (.CLK(net171),
    .D(_0224_),
    .Q(\BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_2 _6210_ (.CLK(net172),
    .D(_0225_),
    .Q(\BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_2 _6211_ (.CLK(net173),
    .D(_0226_),
    .Q(\BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_2 _6212_ (.CLK(net174),
    .D(_0227_),
    .Q(\BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_2 _6213_ (.CLK(net175),
    .D(_0228_),
    .Q(\BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_2 _6214_ (.CLK(net176),
    .D(_0229_),
    .Q(\BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_2 _6215_ (.CLK(net177),
    .D(_0230_),
    .Q(\BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_2 _6216_ (.CLK(net178),
    .D(_0231_),
    .Q(\BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_2 _6217_ (.CLK(net179),
    .D(_0232_),
    .Q(\BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_2 _6218_ (.CLK(net180),
    .D(_0233_),
    .Q(\BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_2 _6219_ (.CLK(net181),
    .D(_0234_),
    .Q(\BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_2 _6220_ (.CLK(net182),
    .D(_0235_),
    .Q(\BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_2 _6221_ (.CLK(net183),
    .D(_0236_),
    .Q(\BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_2 _6222_ (.CLK(net184),
    .D(_0237_),
    .Q(\BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_2 _6223_ (.CLK(net185),
    .D(_0238_),
    .Q(\BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_4 _6224_ (.CLK(net186),
    .D(_0239_),
    .Q(\BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_2 _6225_ (.CLK(net187),
    .D(_0240_),
    .Q(\BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_4 _6226_ (.CLK(net188),
    .D(_0241_),
    .Q(\BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_4 _6227_ (.CLK(net189),
    .D(_0242_),
    .Q(\BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_2 _6228_ (.CLK(net190),
    .D(_0243_),
    .Q(\BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _6229_ (.CLK(net191),
    .D(_0244_),
    .Q(\BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6230_ (.CLK(net192),
    .D(_0245_),
    .Q(\BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6231_ (.CLK(net193),
    .D(_0246_),
    .Q(\BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6232_ (.CLK(net194),
    .D(_0247_),
    .Q(\BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6233_ (.CLK(net195),
    .D(_0248_),
    .Q(\BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6234_ (.CLK(net196),
    .D(_0249_),
    .Q(\BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6235_ (.CLK(net197),
    .D(_0250_),
    .Q(\BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6236_ (.CLK(net38),
    .D(_0251_),
    .Q(\BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6237_ (.CLK(net39),
    .D(_0252_),
    .Q(\BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6238_ (.CLK(net40),
    .D(_0253_),
    .Q(\BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_2 _6239_ (.CLK(net41),
    .D(_0254_),
    .Q(\BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_2 _6240_ (.CLK(net42),
    .D(_0255_),
    .Q(\BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_2 _6241_ (.CLK(net43),
    .D(_0256_),
    .Q(\BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_2 _6242_ (.CLK(net44),
    .D(_0257_),
    .Q(\BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_2 _6243_ (.CLK(net45),
    .D(_0258_),
    .Q(\BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_2 _6244_ (.CLK(net46),
    .D(_0259_),
    .Q(\BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_2 _6245_ (.CLK(net47),
    .D(_0260_),
    .Q(\BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_2 _6246_ (.CLK(net48),
    .D(_0261_),
    .Q(\BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_2 _6247_ (.CLK(net49),
    .D(_0262_),
    .Q(\BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_2 _6248_ (.CLK(net50),
    .D(_0263_),
    .Q(\BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_2 _6249_ (.CLK(net51),
    .D(_0264_),
    .Q(\BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6250_ (.CLK(net52),
    .D(_0265_),
    .Q(\BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _6251_ (.CLK(net53),
    .D(_0266_),
    .Q(\BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _6252_ (.CLK(net54),
    .D(_0267_),
    .Q(\BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_2 _6253_ (.CLK(net55),
    .D(_0268_),
    .Q(\BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_2 _6254_ (.CLK(net56),
    .D(_0269_),
    .Q(\BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_2 _6255_ (.CLK(net57),
    .D(_0270_),
    .Q(\BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_2 _6256_ (.CLK(net58),
    .D(_0271_),
    .Q(\BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_2 _6257_ (.CLK(net59),
    .D(_0272_),
    .Q(\BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_2 _6258_ (.CLK(net60),
    .D(_0273_),
    .Q(\BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_2 _6259_ (.CLK(net61),
    .D(_0274_),
    .Q(\BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_2 _6260_ (.CLK(net62),
    .D(_0275_),
    .Q(\BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_2 _6261_ (.CLK(net63),
    .D(_0276_),
    .Q(\BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_2 _6262_ (.CLK(net64),
    .D(_0277_),
    .Q(\BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_2 _6263_ (.CLK(net65),
    .D(_0278_),
    .Q(\BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_2 _6264_ (.CLK(net66),
    .D(_0279_),
    .Q(\BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_2 _6265_ (.CLK(net67),
    .D(_0280_),
    .Q(\BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_4 _6266_ (.CLK(net68),
    .D(_0281_),
    .Q(\BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_2 _6267_ (.CLK(net69),
    .D(_0282_),
    .Q(\BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6268_ (.CLK(net70),
    .D(_0283_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_2 _6269_ (.CLK(net71),
    .D(_0284_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _6270_ (.CLK(net72),
    .D(_0285_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _6271_ (.CLK(net73),
    .D(_0286_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _6272_ (.CLK(net74),
    .D(_0287_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_2 _6273_ (.CLK(net75),
    .D(_0288_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _6274_ (.CLK(net76),
    .D(_0289_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _6275_ (.CLK(net77),
    .D(_0290_),
    .Q(\BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfxtp_2 _6276_ (.CLK(net78),
    .D(_0291_),
    .Q(\BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6277_ (.CLK(net79),
    .D(_0292_),
    .Q(\BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6278_ (.CLK(net80),
    .D(_0293_),
    .Q(\BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6279_ (.CLK(net81),
    .D(_0294_),
    .Q(\BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6280_ (.CLK(net82),
    .D(_0295_),
    .Q(\BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6281_ (.CLK(net83),
    .D(_0296_),
    .Q(\BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6282_ (.CLK(net84),
    .D(_0297_),
    .Q(\BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6283_ (.CLK(net85),
    .D(_0298_),
    .Q(\BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _6284_ (.CLK(net86),
    .D(_0299_),
    .Q(\BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6285_ (.CLK(net87),
    .D(_0300_),
    .Q(\BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6286_ (.CLK(net88),
    .D(_0301_),
    .Q(\BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6287_ (.CLK(net89),
    .D(_0302_),
    .Q(\BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6288_ (.CLK(net90),
    .D(_0303_),
    .Q(\BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6289_ (.CLK(net91),
    .D(_0304_),
    .Q(\BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6290_ (.CLK(net92),
    .D(_0305_),
    .Q(\BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6291_ (.CLK(net93),
    .D(_0306_),
    .Q(\BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6292_ (.CLK(net94),
    .D(_0307_),
    .Q(\BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6293_ (.CLK(net95),
    .D(_0308_),
    .Q(\BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6294_ (.CLK(net96),
    .D(_0309_),
    .Q(\BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6295_ (.CLK(net97),
    .D(_0310_),
    .Q(\BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6296_ (.CLK(net98),
    .D(_0311_),
    .Q(\BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6297_ (.CLK(net99),
    .D(_0312_),
    .Q(\BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6298_ (.CLK(net100),
    .D(_0313_),
    .Q(\BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6299_ (.CLK(net101),
    .D(_0314_),
    .Q(\BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6300_ (.CLK(net102),
    .D(_0315_),
    .Q(\BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6301_ (.CLK(net103),
    .D(_0316_),
    .Q(\BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _6302_ (.CLK(net104),
    .D(_0317_),
    .Q(\BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6303_ (.CLK(net105),
    .D(_0318_),
    .Q(\BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6304_ (.CLK(net106),
    .D(_0319_),
    .Q(\BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6305_ (.CLK(net107),
    .D(_0320_),
    .Q(\BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6306_ (.CLK(net37),
    .D(_0321_),
    .Q(\BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2580_ (.A(_2580_),
    .X(clknet_0__2580_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2581_ (.A(_2581_),
    .X(clknet_0__2581_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2582_ (.A(_2582_),
    .X(clknet_0__2582_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2583_ (.A(_2583_),
    .X(clknet_0__2583_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2584_ (.A(_2584_),
    .X(clknet_0__2584_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2585_ (.A(_2585_),
    .X(clknet_0__2585_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2586_ (.A(_2586_),
    .X(clknet_0__2586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2587_ (.A(_2587_),
    .X(clknet_0__2587_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2588_ (.A(_2588_),
    .X(clknet_0__2588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2589_ (.A(_2589_),
    .X(clknet_0__2589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2590_ (.A(_2590_),
    .X(clknet_0__2590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2591_ (.A(_2591_),
    .X(clknet_0__2591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2592_ (.A(_2592_),
    .X(clknet_0__2592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2593_ (.A(_2593_),
    .X(clknet_0__2593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2594_ (.A(_2594_),
    .X(clknet_0__2594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2595_ (.A(_2595_),
    .X(clknet_0__2595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2596_ (.A(_2596_),
    .X(clknet_0__2596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2597_ (.A(_2597_),
    .X(clknet_0__2597_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2580_ (.A(clknet_0__2580_),
    .X(clknet_1_0__leaf__2580_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2581_ (.A(clknet_0__2581_),
    .X(clknet_1_0__leaf__2581_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2582_ (.A(clknet_0__2582_),
    .X(clknet_1_0__leaf__2582_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2583_ (.A(clknet_0__2583_),
    .X(clknet_1_0__leaf__2583_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2584_ (.A(clknet_0__2584_),
    .X(clknet_1_0__leaf__2584_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2585_ (.A(clknet_0__2585_),
    .X(clknet_1_0__leaf__2585_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2586_ (.A(clknet_0__2586_),
    .X(clknet_1_0__leaf__2586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2587_ (.A(clknet_0__2587_),
    .X(clknet_1_0__leaf__2587_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2588_ (.A(clknet_0__2588_),
    .X(clknet_1_0__leaf__2588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2589_ (.A(clknet_0__2589_),
    .X(clknet_1_0__leaf__2589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2590_ (.A(clknet_0__2590_),
    .X(clknet_1_0__leaf__2590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2591_ (.A(clknet_0__2591_),
    .X(clknet_1_0__leaf__2591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2592_ (.A(clknet_0__2592_),
    .X(clknet_1_0__leaf__2592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2593_ (.A(clknet_0__2593_),
    .X(clknet_1_0__leaf__2593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2594_ (.A(clknet_0__2594_),
    .X(clknet_1_0__leaf__2594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2595_ (.A(clknet_0__2595_),
    .X(clknet_1_0__leaf__2595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2596_ (.A(clknet_0__2596_),
    .X(clknet_1_0__leaf__2596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2597_ (.A(clknet_0__2597_),
    .X(clknet_1_0__leaf__2597_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2580_ (.A(clknet_0__2580_),
    .X(clknet_1_1__leaf__2580_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2581_ (.A(clknet_0__2581_),
    .X(clknet_1_1__leaf__2581_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2582_ (.A(clknet_0__2582_),
    .X(clknet_1_1__leaf__2582_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2583_ (.A(clknet_0__2583_),
    .X(clknet_1_1__leaf__2583_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2584_ (.A(clknet_0__2584_),
    .X(clknet_1_1__leaf__2584_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2585_ (.A(clknet_0__2585_),
    .X(clknet_1_1__leaf__2585_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2586_ (.A(clknet_0__2586_),
    .X(clknet_1_1__leaf__2586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2587_ (.A(clknet_0__2587_),
    .X(clknet_1_1__leaf__2587_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2588_ (.A(clknet_0__2588_),
    .X(clknet_1_1__leaf__2588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2589_ (.A(clknet_0__2589_),
    .X(clknet_1_1__leaf__2589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2590_ (.A(clknet_0__2590_),
    .X(clknet_1_1__leaf__2590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2591_ (.A(clknet_0__2591_),
    .X(clknet_1_1__leaf__2591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2592_ (.A(clknet_0__2592_),
    .X(clknet_1_1__leaf__2592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2593_ (.A(clknet_0__2593_),
    .X(clknet_1_1__leaf__2593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2594_ (.A(clknet_0__2594_),
    .X(clknet_1_1__leaf__2594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2595_ (.A(clknet_0__2595_),
    .X(clknet_1_1__leaf__2595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2596_ (.A(clknet_0__2596_),
    .X(clknet_1_1__leaf__2596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2597_ (.A(clknet_0__2597_),
    .X(clknet_1_1__leaf__2597_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net30),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_1942_),
    .X(net199));
 sky130_fd_sc_hd__buf_1 hold3 (.A(_1943_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_1944_),
    .X(net201));
 sky130_fd_sc_hd__buf_4 input1 (.A(BitStream_buffer_input[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(BitStream_buffer_input[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(BitStream_buffer_input[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_8 input12 (.A(BitStream_buffer_input[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(BitStream_buffer_input[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(BitStream_buffer_input[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 input15 (.A(BitStream_buffer_input[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(BitStream_buffer_input[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(exp_golomb_sel[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(exp_golomb_sel[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(reset_n),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(BitStream_buffer_input[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(BitStream_buffer_input[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(BitStream_buffer_input[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(BitStream_buffer_input[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(BitStream_buffer_input[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(BitStream_buffer_input[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(BitStream_buffer_input[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(BitStream_buffer_input[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 max_cap35 (.A(_2628_),
    .X(net35));
 sky130_fd_sc_hd__buf_4 max_cap36 (.A(_2620_),
    .X(net36));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(exp_golomb_decoding_output[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(exp_golomb_decoding_output[1]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(exp_golomb_decoding_output[2]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(exp_golomb_decoding_output[3]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(exp_golomb_decoding_output[4]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(exp_golomb_decoding_output[5]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(exp_golomb_decoding_output[6]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(exp_golomb_decoding_output[7]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(half_fill_counter[0]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(half_fill_counter[1]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(half_fill_counter[2]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(reset_counter[0]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(reset_counter[1]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(reset_counter[2]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(reset_counter[3]));
endmodule

