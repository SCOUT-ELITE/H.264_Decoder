* NGSPICE file created from egd_top_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

.subckt egd_top_wrapper la_data_in_47_32[0] la_data_in_47_32[10] la_data_in_47_32[11]
+ la_data_in_47_32[12] la_data_in_47_32[13] la_data_in_47_32[14] la_data_in_47_32[15]
+ la_data_in_47_32[1] la_data_in_47_32[2] la_data_in_47_32[3] la_data_in_47_32[4]
+ la_data_in_47_32[5] la_data_in_47_32[6] la_data_in_47_32[7] la_data_in_47_32[8]
+ la_data_in_47_32[9] la_data_in_49_48[0] la_data_in_49_48[1] la_data_in_65 la_data_out_15_8[0]
+ la_data_out_15_8[1] la_data_out_15_8[2] la_data_out_15_8[3] la_data_out_15_8[4]
+ la_data_out_15_8[5] la_data_out_15_8[6] la_data_out_15_8[7] la_data_out_18_16[0]
+ la_data_out_18_16[1] la_data_out_18_16[2] la_data_out_22_19[0] la_data_out_22_19[1]
+ la_data_out_22_19[2] la_data_out_22_19[3] vccd1 vssd1 wb_clk_i
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3988_ _3108_ _3077_ _0703_ _0704_ _0705_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5727_ net15 _3105_ _2353_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5658_ _2324_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4609_ _0923_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _1323_
+ sky130_fd_sc_hd__or2b_1
X_5589_ net16 _0469_ _2281_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6217__84 clknet_1_0__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
XFILLER_0_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4960_ _0574_ _0963_ _3075_ _0964_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4891_ _2800_ _0787_ _3097_ _0788_ _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3911_ _2870_ _2872_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3842_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__inv_2
X_5512_ _0885_ _0414_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__nand2_1
X_3773_ _0392_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6492_ net66 egd_top.BitStream_buffer.pc\[0\] net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5443_ _0920_ _0945_ _0946_ _0346_ _2149_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__a221oi_1
X_5374_ _2887_ _0840_ _3010_ _0842_ _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__a221oi_1
X_4325_ _0926_ _0831_ _0832_ _2816_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4256_ _0967_ _0625_ _0968_ _0777_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__a221oi_1
X_3207_ _2773_ _2774_ _2775_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__and3_1
X_4187_ _0385_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2722_ clknet_0__2722_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2722_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4110_ _3012_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__clkbuf_4
X_5090_ _2848_ _0996_ _0495_ _0997_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4041_ _0411_ _2887_ _0413_ _3007_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5992_ _2505_ _2439_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4943_ _1640_ _1644_ _1649_ _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4874_ _0941_ _0709_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3825_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3756_ _2896_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0475_
+ sky130_fd_sc_hd__nand2_1
X_6475_ net217 _0308_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[124\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3687_ _0406_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
X_5426_ _3122_ _2931_ _3125_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1
+ vccd1 vccd1 _2133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5357_ _2053_ _2056_ _2059_ _2063_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__and4_2
X_4308_ _0802_ _0330_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__nand2_1
X_5288_ _0981_ _2920_ _0982_ _2922_ _1995_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__a221oi_1
X_4239_ _3152_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3610_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _0895_ _2828_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__nand2_1
X_3541_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3472_ _3020_ _2808_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5211_ _3034_ _0922_ _2904_ _0921_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__a221oi_1
X_5142_ _1840_ _1844_ _1846_ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__and4_1
X_5073_ _2818_ _0954_ _2816_ _0955_ _1782_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__a221oi_2
X_4024_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__clkbuf_8
X_6265__128 clknet_1_1__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5975_ _2551_ _2512_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4926_ _0865_ _3132_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2724_ _2724_ vssd1 vssd1 vccd1 vccd1 clknet_0__2724_ sky130_fd_sc_hd__clkbuf_16
X_4857_ _2887_ _0987_ _2881_ _0989_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ _3033_ _3048_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nand2_1
X_4788_ _0820_ _2820_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__nand2_1
X_3739_ _0458_ _0456_ _2789_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__o21ai_1
X_6458_ net200 _0291_ net38 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5409_ _0999_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _2116_
+ sky130_fd_sc_hd__nand2_1
X_6389_ net131 _0222_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6187__56 clknet_1_0__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__inv_2
XFILLER_0_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5760_ net5 _0443_ _2377_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5691_ net16 egd_top.BitStream_buffer.BS_buffer\[54\] _2335_ vssd1 vssd1 vccd1 vccd1
+ _2342_ sky130_fd_sc_hd__mux2_1
X_4711_ _1410_ _1414_ _1419_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4642_ _1354_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__nand2_1
X_4573_ _0341_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__inv_2
X_3524_ _3042_ _3052_ _3063_ _3072_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__and4_1
X_3455_ _2895_ _2961_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__and2_1
X_3386_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__buf_6
X_5125_ _0804_ _1011_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5056_ _0984_ _0882_ _1763_ _1764_ _1765_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__o2111a_1
X_4007_ _2802_ _3157_ _0329_ _2800_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5958_ _2500_ _2534_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__nand2_1
X_4909_ _0833_ _2820_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5889_ _2464_ _2465_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6248__112 clknet_1_1__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_5 _0505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3240_ net5 _2802_ _2798_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__mux2_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _2740_ _2741_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__nor2_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5812_ _2412_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5743_ net1 _2959_ _2352_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5674_ _2332_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4625_ _3031_ _0956_ _0698_ _0958_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__o22ai_1
X_4556_ _0816_ _3066_ _0817_ _2824_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__a221oi_1
X_3507_ _2933_ _2996_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4487_ _0881_ _3080_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__or2_1
X_3438_ egd_top.BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__clkbuf_8
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _2908_ _2912_ _2914_ _2917_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__o22ai_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _1816_ _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__nor2_1
X_6088_ _2656_ _2657_ _2513_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__o21ai_1
X_5039_ _2935_ _0857_ _0378_ _0858_ _1748_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[0] sky130_fd_sc_hd__buf_12
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[0] sky130_fd_sc_hd__buf_12
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__clkinv_4
X_5390_ _2095_ _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__nand2_1
X_4341_ _0867_ _3119_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nand2_1
X_4272_ _0417_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__buf_4
X_6011_ _2581_ _2586_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__nor2_1
X_3223_ net221 vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__inv_2
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3987_ _3087_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0705_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5726_ _2360_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5657_ net16 _0341_ _2317_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5588_ _2287_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__clkbuf_1
X_4608_ _1311_ _1314_ _1317_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__and4_1
X_4539_ _0791_ _2990_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4890_ _0957_ _0790_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__o21ai_1
X_3910_ _0627_ _0628_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__nand2_1
X_3841_ _3123_ _0395_ _3126_ _3124_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3772_ _2949_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _0491_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5511_ _0883_ _2887_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6491_ net65 _0324_ net35 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5442_ _2147_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__nand2_1
X_5373_ _0407_ _0843_ _2079_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__o21ai_1
X_4324_ _1038_ _1039_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _3075_ _0969_ _0970_ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__o22ai_1
X_3206_ egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 _2775_
+ sky130_fd_sc_hd__inv_2
X_4186_ _0456_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5709_ net1 _3142_ _2334_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__2721_ clknet_0__2721_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2721_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _0756_ _0405_ _0757_ _0409_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5991_ _2481_ _2499_ _2443_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4942_ _0892_ _2848_ _0893_ _0587_ _1652_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4873_ _0939_ _0336_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3824_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3755_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3686_ egd_top.BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6474_ net216 _0307_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[125\]
+ sky130_fd_sc_hd__dfrtp_4
X_5425_ _1185_ _3076_ _2129_ _2130_ _2131_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5356_ _2810_ _0800_ _0801_ _0625_ _2062_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4307_ _1021_ _3065_ _0957_ _0796_ _1022_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__o221a_1
X_5287_ _1052_ _0404_ _2908_ _0408_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__o22ai_1
X_4238_ _0329_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__buf_8
X_4169_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__clkbuf_8
X_6242__107 clknet_1_1__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3540_ _3075_ _3077_ _3081_ _3085_ _3088_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5210_ _0465_ _0923_ _1918_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__o21ai_1
X_3471_ _2870_ _2996_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__and2_1
X_5141_ _0420_ _0831_ _0832_ _0458_ _1849_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__a221oi_1
X_5072_ _1017_ _0956_ _1256_ _0958_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ _2957_ _0368_ _0370_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1
+ vccd1 vccd1 _0741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5974_ _2528_ _2550_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4925_ _1627_ _1630_ _1633_ _1635_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4856_ _1566_ _1567_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__2723_ _2723_ vssd1 vssd1 vccd1 vccd1 clknet_0__2723_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3807_ _3037_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__clkinv_4
X_4787_ _0818_ _2826_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3738_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3669_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__buf_4
X_6457_ net199 _0290_ net38 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_5408_ _0427_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _2115_
+ sky130_fd_sc_hd__nand2_1
X_6388_ net130 _0221_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[68\]
+ sky130_fd_sc_hd__dfrtp_2
X_5339_ _2023_ _2037_ _2046_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5690_ _2341_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4710_ _0892_ _2830_ _0893_ _0920_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4641_ _0999_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _1355_
+ sky130_fd_sc_hd__nand2_1
X_4572_ _0657_ _2840_ _2847_ _1000_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__a221oi_1
X_3523_ _3064_ _3065_ _3067_ _3068_ _3071_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__o221a_1
X_3454_ _3001_ _3002_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__nand2_1
X_6271__133 clknet_1_0__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
X_3385_ _2933_ _2910_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__and2_1
X_5124_ _0802_ _2810_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__nand2_1
X_5055_ _0889_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _1765_
+ sky130_fd_sc_hd__or2b_1
X_4006_ _0619_ _3152_ _0723_ _3155_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5957_ _2532_ _2533_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4908_ _0824_ _3090_ _0825_ _2907_ _1618_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5888_ egd_top.BitStream_buffer.BitStream_buffer_valid_n egd_top.BitStream_buffer.BitStream_buffer_output\[15\]
+ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__nor2_1
X_4839_ _3008_ _3084_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 _0546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6294__155 clknet_1_1__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__inv_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ net31 _2737_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5811_ net36 egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__nand2_1
X_6314__5 clknet_1_1__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__inv_2
XFILLER_0_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5742_ _2368_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5673_ net8 egd_top.BitStream_buffer.BS_buffer\[46\] _2316_ vssd1 vssd1 vccd1 vccd1
+ _2332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4624_ _1326_ _1329_ _1333_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__and4_1
X_4555_ _1267_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__nand2_1
X_6323__13 clknet_1_0__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__inv_2
XFILLER_0_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3506_ _3054_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__buf_1
X_4486_ _0395_ _3096_ _3104_ _0463_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__a221oi_1
X_3437_ _2895_ _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__and2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _2916_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__clkbuf_4
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5107_ _0933_ _0638_ _0934_ _0610_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__a22o_1
X_6087_ _2655_ _2650_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__and2_1
X_3299_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__clkbuf_8
X_5038_ _3144_ _2912_ _1287_ _2917_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[1] sky130_fd_sc_hd__buf_12
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[1] sky130_fd_sc_hd__buf_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6302__162 clknet_1_0__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__inv_2
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6171__41 clknet_1_0__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__inv_2
XFILLER_0_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4340_ _0865_ _2974_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__nand2_1
X_4271_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__buf_6
X_3222_ _2788_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__clkbuf_1
X_6010_ _2582_ _2583_ _2496_ _2585_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__2729_ clknet_0__2729_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2729_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3986_ _3078_ _3084_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5725_ net16 _0656_ _2353_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5656_ _2323_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4607_ _0904_ _3077_ _1318_ _1319_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__o2111a_1
X_5587_ net2 _2874_ _2281_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__mux2_1
X_4538_ _1011_ _0781_ _3058_ _0782_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4469_ _0885_ _0469_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__nand2_1
X_6139_ _2705_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__inv_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6208__75 clknet_1_0__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3840_ _3129_ _3110_ _0556_ _0557_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6223__89 clknet_1_0__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
XFILLER_0_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3771_ _2947_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _0490_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5510_ _0892_ _0894_ _0893_ _0607_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6490_ net64 _0323_ net36 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ _0949_ _0553_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__nand2_1
X_5372_ _0844_ _3058_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__nand2_1
X_4323_ _0835_ _2826_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4254_ _0350_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3205_ egd_top.BitStream_buffer.buffer_index\[5\] vssd1 vssd1 vccd1 vccd1 _2774_
+ sky130_fd_sc_hd__inv_2
X_4185_ _0808_ _0839_ _0862_ _0901_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3969_ _3033_ _3002_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__nand2_1
X_5708_ _2350_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5639_ net8 _3097_ _2298_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__2720_ clknet_0__2720_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2720_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _2508_ _2522_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4941_ _1650_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4872_ _0657_ _0945_ _0946_ _3132_ _1583_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3823_ _0484_ _0505_ _0525_ _0541_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__and4_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3754_ _2920_ _2867_ _2873_ _0469_ _0472_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__a221oi_1
X_3685_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6473_ net215 _0306_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[126\]
+ sky130_fd_sc_hd__dfrtp_4
X_5424_ _3086_ _0435_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5355_ _2060_ _2061_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4306_ _0797_ _2802_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__nand2_1
X_5286_ _1950_ _1964_ _1976_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__and4_1
X_4237_ _3157_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__buf_6
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4168_ _2949_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__clkbuf_4
X_4099_ _3001_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3470_ _3013_ _3018_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__nor2_1
X_5140_ _1847_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__nand2_1
X_5071_ _1770_ _1773_ _1776_ _1780_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__and4_1
X_4022_ _0736_ _0737_ _0738_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5973_ _2536_ _2549_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__nor2_1
X_4924_ _0395_ _0857_ _2935_ _0858_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_19_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2722_ _2722_ vssd1 vssd1 vccd1 vccd1 clknet_0__2722_ sky130_fd_sc_hd__clkbuf_16
X_4855_ _0992_ _3037_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4786_ _2802_ _0810_ _3058_ _0809_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__a221oi_1
X_3806_ _0510_ _0515_ _0519_ _0524_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__and4_1
X_3737_ _0456_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__clkbuf_4
X_3668_ _2878_ _2937_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__and2_1
X_6456_ net198 _0289_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3599_ _2878_ _2910_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__nand2_1
X_5407_ _3040_ _0987_ _3007_ _0989_ _2113_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__a221oi_1
X_6387_ net129 _0220_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[69\]
+ sky130_fd_sc_hd__dfrtp_2
X_5338_ _2039_ _2041_ _2043_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__and4_2
X_5269_ _0865_ _2939_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4640_ _0428_ _0894_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4571_ _1005_ _2854_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__o21ai_1
X_3522_ _3069_ _3070_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3453_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__buf_4
X_5123_ _2822_ _2996_ _2927_ _1831_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__a31oi_1
X_3384_ _2932_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__clkbuf_4
X_5054_ _0885_ _0551_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__nand2_1
X_4005_ _0330_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5956_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__nand2_1
X_4907_ _0756_ _0826_ _2914_ _0827_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__o22ai_1
X_5887_ _2462_ _2463_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4838_ _3011_ _3080_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4769_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] vssd1 vssd1 vccd1
+ vccd1 _1482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6439_ net181 _0272_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_7 _0546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5810_ _2411_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[4\] sky130_fd_sc_hd__buf_2
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5741_ net8 _0464_ _2352_ vssd1 vssd1 vccd1 vccd1 _2368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5672_ _2331_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4623_ _2959_ _0945_ _0946_ _0336_ _1336_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4554_ _0820_ _2816_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3505_ _2864_ _2984_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4485_ _1052_ _3093_ _1199_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__o21ai_1
X_3436_ _2984_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__buf_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _2878_ _2915_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__nand2_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ egd_top.BitStream_buffer.BS_buffer\[76\] _0930_ _0931_ egd_top.BitStream_buffer.BS_buffer\[79\]
+ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a22o_1
X_6086_ _2650_ _2655_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__nor2_2
X_3298_ _2846_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__buf_4
X_5037_ _0926_ _2840_ _2847_ _0875_ _1746_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6229__95 clknet_1_1__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5939_ _2515_ _2482_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__nand2_2
X_6157__28 clknet_1_0__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__inv_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[2] sky130_fd_sc_hd__buf_12
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[2] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ _0422_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__buf_4
X_3221_ _2787_ net28 _2783_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2728_ clknet_0__2728_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2728_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3985_ _2944_ _3080_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5724_ _2359_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
X_5655_ net2 _0378_ _2317_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4606_ _3087_ _0389_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__nand2_1
X_5586_ _2286_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__clkbuf_1
X_4537_ egd_top.BitStream_buffer.BS_buffer\[1\] _0783_ _0784_ _0777_ vssd1 vssd1 vccd1
+ vccd1 _1251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4468_ _0883_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _1183_
+ sky130_fd_sc_hd__nand2_1
X_3419_ _2956_ _2957_ _2958_ _2959_ _2967_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__a221oi_1
X_6138_ _2704_ _2512_ _2505_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__nand3_1
X_4399_ _0981_ _2993_ _0982_ _3010_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__a221oi_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _2636_ _2638_ _2509_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3770_ _0412_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5440_ _0947_ _0656_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5371_ _2067_ _2071_ _2073_ _2077_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ _0833_ _2810_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4253_ _2926_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__inv_2
X_3204_ egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 _2773_
+ sky130_fd_sc_hd__inv_2
X_4184_ _0870_ _0880_ _0891_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3968_ _3053_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__clkinv_4
X_5707_ net8 _0392_ _2334_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3899_ _0439_ egd_top.BitStream_buffer.BS_buffer\[91\] _0441_ egd_top.BitStream_buffer.BS_buffer\[92\]
+ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5638_ _2313_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5569_ _2251_ _2265_ _2274_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4940_ _0897_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _1651_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4871_ _1581_ _1582_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3822_ _0530_ _0533_ _0537_ _0540_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3753_ _0470_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3684_ _2964_ _2915_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6472_ net214 _0305_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[127\]
+ sky130_fd_sc_hd__dfrtp_4
X_5423_ _0757_ _3083_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5354_ _0804_ _2874_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__nand2_1
X_4305_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5285_ _1980_ _1984_ _1988_ _1992_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__and4_1
X_4236_ _0929_ _0936_ _0944_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__and4_2
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _0883_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _0884_
+ sky130_fd_sc_hd__nand2_1
X_4098_ _3002_ _0809_ _3153_ _0810_ _0814_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6199__67 clknet_1_1__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__inv_2
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _0653_ _3077_ _1777_ _1778_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__o2111a_1
X_4021_ _0363_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _0739_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5972_ _2540_ _2548_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4923_ _0334_ _2912_ _1171_ _2917_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_0__2721_ _2721_ vssd1 vssd1 vccd1 vccd1 clknet_0__2721_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4854_ _0990_ _3034_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4785_ _1171_ _0811_ _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3805_ _0520_ _0521_ _0522_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3736_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__buf_2
X_3667_ _0379_ _0381_ _0383_ _0386_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6455_ net197 _0288_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3598_ _3146_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__inv_2
X_6386_ net128 _0219_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[70\]
+ sky130_fd_sc_hd__dfrtp_2
X_5406_ _2111_ _2112_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5337_ _0974_ _0346_ _0975_ _3112_ _2044_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__a221oi_1
X_5268_ _1967_ _1970_ _1973_ _1975_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__and4_1
X_4219_ _0932_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nor2_1
X_5199_ _1906_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6178__48 clknet_1_1__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__inv_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4570_ _2858_ _0495_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3521_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3452_ _2899_ _2985_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3383_ _2876_ egd_top.BitStream_buffer.pc\[2\] _2868_ vssd1 vssd1 vccd1 vccd1 _2932_
+ sky130_fd_sc_hd__and3_1
X_5122_ _1256_ _0796_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5053_ _0883_ _2881_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__nand2_1
X_4004_ _0366_ _3141_ _2771_ _0398_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5955_ _2531_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _0816_ _0330_ _0817_ _0458_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5886_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] egd_top.BitStream_buffer.BitStream_buffer_output\[14\]
+ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4837_ _0341_ _3096_ _3104_ _2959_ _1548_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4768_ _1479_ _1480_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4699_ _0877_ _2931_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__nand2_1
X_6438_ net180 _0271_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6369_ net111 _0202_ net42 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 _0755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6255__119 clknet_1_0__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5740_ _2367_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5671_ net9 _3132_ _2316_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__mux2_1
X_4622_ _1334_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__nand2_1
X_4553_ _0818_ _2822_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3504_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__clkbuf_8
X_4484_ _3100_ _0414_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3435_ _2983_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__inv_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _2865_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__clkbuf_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _0937_ _0656_ _0553_ _0938_ _1814_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__a221oi_1
X_6085_ _2654_ _2619_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__nand2_1
X_3297_ _2845_ _2837_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__and2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5036_ _0686_ _2854_ _1745_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5938_ _2499_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5869_ _2444_ _2445_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[3] sky130_fd_sc_hd__buf_12
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[3] sky130_fd_sc_hd__buf_12
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3220_ net28 _2752_ _2778_ _2780_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2727_ clknet_0__2727_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2727_
+ sky130_fd_sc_hd__clkbuf_16
X_3984_ _0645_ _0667_ _0685_ _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5723_ net2 _0371_ _2353_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5654_ _2322_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4605_ _0650_ _3084_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__or2_1
X_6238__103 clknet_1_0__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5585_ net3 _0886_ _2281_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4536_ _1249_ _1250_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4467_ _0607_ _0872_ _1000_ _0873_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__a221oi_1
X_4398_ _2914_ _0405_ _0403_ _0409_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o22ai_1
X_3418_ _2963_ _2966_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__nand2_1
X_6137_ _2684_ _2683_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__or2_1
X_3349_ _2855_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__inv_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _2637_ _2634_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__nand2_1
X_5019_ _0820_ _2824_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__nand2_1
X_6284__145 clknet_1_1__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
XFILLER_0_67_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5370_ _2904_ _0831_ _0832_ _0777_ _2076_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__a221oi_1
X_4321_ _0824_ _2920_ _0825_ _2922_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__a221oi_1
X_4252_ _0348_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__clkbuf_4
X_3203_ _2753_ _2757_ egd_top.BitStream_buffer.pc\[6\] _2771_ vssd1 vssd1 vccd1 vccd1
+ _2772_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4183_ _0892_ _3105_ _0893_ _0894_ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3967_ _0671_ _0676_ _0679_ _0684_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5706_ _2349_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3898_ _0613_ _0614_ _0615_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__and4_1
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5637_ net9 _2980_ _2298_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5568_ _2267_ _2269_ _2271_ _2273_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4519_ _0990_ _0610_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__nand2_1
X_5499_ _0865_ _0346_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__nand2_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6213__80 clknet_1_1__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4870_ _0949_ _0435_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3821_ _0538_ _3065_ _3154_ _3068_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3752_ _2886_ _3007_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3683_ _0402_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
X_6471_ net213 _0304_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_5422_ _0403_ _3079_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__or2_1
X_5353_ _0802_ _2814_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__nand2_1
X_4304_ _3066_ _0787_ _2863_ _0788_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _0601_ _0882_ _1989_ _1990_ _1991_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__o2111a_1
X_4235_ _0463_ _0945_ _0946_ _2974_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4166_ _2947_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__clkbuf_4
X_4097_ _2908_ _0811_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4999_ _1708_ _1709_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4020_ _0361_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0738_
+ sky130_fd_sc_hd__nand2_1
X_5971_ _2547_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4922_ _0830_ _2840_ _2847_ _0920_ _1632_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__a221oi_1
Xclkbuf_0__2720_ _2720_ vssd1 vssd1 vccd1 vccd1 clknet_0__2720_ sky130_fd_sc_hd__clkbuf_16
X_4853_ _0981_ _3015_ _0982_ _3017_ _1564_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4784_ _0812_ _2920_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3804_ _3026_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _0523_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3735_ egd_top.BitStream_buffer.pc\[6\] egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\]
+ _0454_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6454_ net196 _0287_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3666_ _0384_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__nand2_1
X_5405_ _0992_ _3153_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6385_ net127 _0218_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[71\]
+ sky130_fd_sc_hd__dfrtp_4
X_3597_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__clkbuf_8
X_5336_ _3075_ _0976_ _3108_ _0977_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__o22ai_1
X_5267_ _0341_ _0857_ _0343_ _0858_ _1974_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__a221oi_1
X_4218_ _0933_ _0742_ _0934_ _0583_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__a22o_1
X_5198_ _0992_ _3058_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__nand2_1
X_4149_ _0865_ _0343_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3520_ _2902_ _2985_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3451_ _2999_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _3000_
+ sky130_fd_sc_hd__nand2_1
X_3382_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__buf_4
X_5121_ _0797_ _2816_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__nand2_1
X_5052_ _0892_ _0464_ _0893_ _0742_ _1761_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__a221oi_1
X_4003_ _3147_ _3145_ _0349_ _3148_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5954_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4905_ _1614_ _1615_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__nand2_1
X_5885_ _2460_ _2461_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4836_ _1403_ _3093_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4767_ _0988_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3718_ _2856_ _2851_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__and2_1
X_4698_ _0874_ _0871_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nand2_1
X_6437_ net179 _0270_ net41 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_3649_ _2870_ _2836_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nand2_1
X_6368_ net110 _0201_ net42 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5319_ _3151_ _0923_ _2026_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _0757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6183__52 clknet_1_1__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__inv_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5670_ _2330_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _0949_ _0398_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__nand2_1
X_4552_ _2791_ _0810_ _3053_ _0809_ _1265_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3503_ _3045_ _3051_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__nor2_1
X_4483_ egd_top.BitStream_buffer.BS_buffer\[56\] _0907_ _3142_ _0908_ _1197_ vssd1
+ vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3434_ egd_top.BitStream_buffer.pc\[4\] _2768_ _2835_ vssd1 vssd1 vccd1 vccd1 _2983_
+ sky130_fd_sc_hd__or3_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6153_ clknet_1_1__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__buf_1
X_3365_ _2913_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__inv_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _2551_ _2588_ _2615_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__o21bai_1
X_5104_ _1812_ _1813_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__nand2_1
X_3296_ _2844_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__buf_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _2858_ _0830_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5937_ _2513_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5868_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1 vccd1
+ _2445_ sky130_fd_sc_hd__inv_2
X_5799_ _2404_ egd_top.BitStream_buffer.pc_reg\[4\] vssd1 vssd1 vccd1 vccd1 _2405_
+ sky130_fd_sc_hd__nand2_1
X_4819_ _0883_ _3101_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[4] sky130_fd_sc_hd__buf_12
XFILLER_0_31_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6261__124 clknet_1_1__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_0_39_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2726_ clknet_0__2726_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2726_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5722_ _2358_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__clkbuf_1
X_3983_ _0690_ _0693_ _0697_ _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5653_ net3 _2935_ _2317_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5584_ _2285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__clkbuf_1
X_4604_ _3008_ _3080_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4535_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] vssd1 vssd1
+ vccd1 vccd1 _1250_ sky130_fd_sc_hd__nand2_1
X_6162__33 clknet_1_1__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__inv_2
XFILLER_0_40_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4466_ _1179_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__nand2_1
X_4397_ _1106_ _1108_ _1110_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6205_ clknet_1_1__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__buf_1
X_3417_ _2965_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _2966_
+ sky130_fd_sc_hd__nand2_1
X_6136_ _2701_ _2703_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__nand2_1
X_3348_ _2896_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _2897_
+ sky130_fd_sc_hd__nand2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _2566_ _2631_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__nor2_1
X_3279_ net1 _2828_ _2797_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__mux2_1
X_5018_ _0818_ _0458_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4320_ _0602_ _0826_ _0984_ _0827_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_10_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4251_ _0353_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3202_ _2770_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__buf_6
X_4182_ _0896_ _0898_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3966_ _0680_ _0681_ _0682_ _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__and4_1
X_5705_ net9 _2951_ _2334_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5636_ _2312_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
X_3897_ _0434_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _0616_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5567_ _0974_ _3119_ _0975_ egd_top.BitStream_buffer.BS_buffer\[53\] _2272_ vssd1
+ vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4518_ _0981_ _3010_ _0982_ _0406_ _1232_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__a221oi_1
X_5498_ _2195_ _2198_ _2201_ _2203_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__and4_1
X_4449_ _1116_ _0840_ _0551_ _0842_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__a221oi_1
X_6119_ _2637_ _2682_ _2684_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__nand3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6267__130 clknet_1_0__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3820_ _3069_ _0330_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3751_ _2880_ _2943_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3682_ egd_top.BitStream_buffer.BS_buffer\[24\] vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__buf_4
X_6470_ net212 _0303_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5421_ _0336_ _3095_ _3103_ egd_top.BitStream_buffer.BS_buffer\[84\] _2127_ vssd1
+ vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__a221oi_2
X_5352_ _2826_ _2996_ _2927_ _2058_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__a31oi_1
X_4303_ _1017_ _0790_ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5283_ _0889_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _1991_
+ sky130_fd_sc_hd__or2b_1
X_4234_ _0948_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4165_ _2945_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__buf_4
X_4096_ _0812_ _3040_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nand2_1
X_4998_ _0841_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__o21a_1
X_3949_ _0649_ _0655_ _0661_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5619_ net3 _0406_ _2299_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6317__8 clknet_1_0__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__inv_2
X_5970_ _2541_ _2494_ _2546_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__o21ai_1
X_4921_ _0526_ _2854_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__o21ai_1
X_4852_ _2908_ _0405_ _2914_ _0409_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__o22ai_1
X_3803_ _3024_ _2804_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nand2_1
X_4783_ _1484_ _1487_ _1490_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3734_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] egd_top.BitStream_buffer.pc\[1\]
+ egd_top.BitStream_buffer.pc\[0\] _2872_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__o41a_1
X_3665_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__buf_4
X_6453_ net195 _0286_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5404_ _0990_ _3053_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3596_ _2856_ _2910_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__nand2_1
X_6384_ net126 _0217_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5335_ _0967_ _3101_ _0968_ _0551_ _2042_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__a221oi_1
X_5266_ _3147_ _2911_ _1519_ _2916_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _0374_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__clkbuf_4
X_5197_ _0990_ _3030_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__nand2_1
X_4148_ _2934_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _3068_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3450_ _2899_ _2996_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3381_ _2767_ _2910_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__and2_2
X_5120_ _2804_ _0787_ _2907_ _0788_ _1828_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__a221oi_1
X_5051_ _1759_ _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__nand2_1
X_4002_ _0706_ _0711_ _0715_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5953_ _2501_ _2529_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__nand2_1
X_4904_ _0820_ _2822_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5884_ _2453_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__a21oi_1
X_6169__39 clknet_1_1__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__inv_2
X_4835_ _3100_ _2993_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4766_ _1425_ _0903_ _1478_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3717_ _0429_ _0431_ _0433_ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4697_ egd_top.BitStream_buffer.BS_buffer\[56\] _0863_ _0864_ egd_top.BitStream_buffer.BS_buffer\[54\]
+ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__a221oi_2
X_6436_ net178 _0269_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_3648_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
X_3579_ _3123_ _3124_ _3126_ _3127_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__a22o_1
X_6367_ net109 _0200_ net42 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5318_ _0925_ _2904_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__nand2_1
X_5249_ _0816_ _2802_ _0817_ _1011_ _1956_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_38_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _0947_ _3142_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4551_ _0859_ _0811_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4482_ _1075_ _3110_ _1196_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3502_ _3047_ _3048_ egd_top.BitStream_buffer.BS_buffer\[125\] _3050_ vssd1 vssd1
+ vccd1 vccd1 _3051_ sky130_fd_sc_hd__a22o_1
X_3433_ _2845_ _2915_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__nand2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__clkbuf_8
X_5103_ _0941_ _2830_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _2649_ _2652_ _2514_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__o21ai_1
X_3295_ _2843_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__and3_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _3015_ _0848_ _2920_ _0849_ _1743_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5936_ _2511_ _2512_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5867_ _2442_ _2443_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5798_ _2401_ _2402_ _2403_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__a21bo_1
X_4818_ _0638_ _0872_ _0920_ _0873_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4749_ _0974_ _3132_ _0975_ egd_top.BitStream_buffer.BS_buffer\[46\] _1461_ vssd1
+ vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6419_ net161 _0252_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[37\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[5] sky130_fd_sc_hd__buf_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3982_ _0698_ _3065_ _0567_ _3068_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0__f__2725_ clknet_0__2725_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2725_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ net3 _2957_ _2353_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5652_ _2321_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
X_5583_ net4 _1011_ _2281_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__mux2_1
X_4603_ _2935_ _3096_ _3104_ _2848_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4534_ _1247_ _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4465_ _0877_ _3132_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__nand2_1
X_4396_ _0974_ _3143_ _0975_ _0336_ _1111_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__a221oi_1
X_3416_ _2964_ _2837_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__and2_1
X_6135_ _2677_ _2702_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__nand2_1
X_3347_ _2895_ _2872_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__and2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _2566_ _2631_ _2635_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__o21ai_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5017_ _2806_ _0810_ _3153_ _0809_ _1726_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__a221oi_1
X_3278_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__buf_4
X_6245__109 clknet_1_1__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5919_ _2495_ _2466_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _0352_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__clkbuf_4
X_3201_ _2767_ _2769_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__and2_1
X_4181_ _0897_ _2830_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ _3026_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _0683_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5704_ _2348_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
X_3896_ _0432_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _0615_
+ sky130_fd_sc_hd__nand2_1
X_5635_ net10 _2913_ _2298_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5566_ _3108_ _0976_ _0561_ _0977_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4517_ _2981_ _0405_ _0601_ _0409_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__o22ai_1
X_5497_ _2974_ _0857_ _0333_ _0858_ _2202_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__a221oi_1
X_6290__151 clknet_1_0__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__inv_2
X_4448_ _0544_ _0843_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__o21ai_1
X_4379_ _1093_ _1094_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nor2_1
X_6118_ _2683_ _2685_ vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ net20 net21 vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3750_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__clkbuf_8
X_3681_ _0365_ _0376_ _0387_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__and4_1
X_5420_ _3147_ _3092_ _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__o21ai_1
X_5351_ _1488_ _0796_ _2057_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__o21ai_1
X_4302_ _0791_ _3037_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5282_ _0885_ _2943_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__nand2_1
X_4233_ _0949_ _0392_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nand2_1
X_4164_ _2887_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__inv_2
X_4095_ _2992_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _1655_ _0903_ _1707_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3948_ _0662_ _0663_ _0664_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3879_ _0397_ _0366_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5618_ _2303_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__clkbuf_1
X_5549_ _0619_ _0923_ _2254_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6297__157 clknet_1_0__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__inv_2
XFILLER_0_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4920_ _2858_ _1000_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__nand2_1
X_4851_ _1556_ _1558_ _1560_ _1562_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3802_ _3022_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0521_
+ sky130_fd_sc_hd__nand2_1
X_4782_ _2800_ _0800_ _0801_ _2822_ _1493_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__a221oi_1
X_3733_ _3138_ _0356_ _0401_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3664_ _2833_ _2937_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__and2_1
X_6452_ net194 _0285_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_5403_ _0981_ _2922_ _0982_ _2913_ _2109_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3595_ _3143_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__inv_2
X_6383_ net125 _0216_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[73\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5334_ _0492_ _0969_ _0717_ _0971_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__o22ai_1
X_5265_ _0875_ _2840_ _2847_ _0742_ _1972_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__a221oi_1
X_4216_ _0373_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__clkbuf_4
X_5196_ _0981_ _2863_ _0982_ _2920_ _1904_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4147_ _2930_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__buf_4
X_4078_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3380_ _2928_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__clkbuf_2
X_5050_ _0897_ _0894_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__nand2_1
X_4001_ _0716_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5952_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4903_ _0818_ _2828_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5883_ _2452_ _2459_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__nand2_1
X_4834_ _0385_ _0907_ _0366_ _0908_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4765_ _1438_ _1454_ _1463_ _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3716_ _0434_ _0435_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4696_ _1407_ _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ net177 _0268_ net41 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3647_ _2946_ _2836_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__nand2_1
X_6366_ net108 _0199_ net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_3578_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__clkbuf_8
X_5317_ _0443_ _0933_ _2987_ _0934_ _2024_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__a221oi_1
X_5248_ _1954_ _1955_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__nand2_1
X_5179_ _3144_ _3093_ _1887_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4550_ _0812_ _0402_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__nand2_1
X_3501_ _3049_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__inv_2
X_4481_ _3118_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _1196_
+ sky130_fd_sc_hd__nand2_1
X_3432_ _2980_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__inv_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _2562_ _2513_ _2554_ _2716_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__a31o_1
X_3363_ _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__clkbuf_4
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _0939_ _3132_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__nand2_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _2650_ _2651_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__nor2_1
X_3294_ _2842_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__inv_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _0650_ _0850_ _1742_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5935_ _2760_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5866_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1 vccd1
+ _2443_ sky130_fd_sc_hd__inv_2
X_4817_ _1527_ _1528_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5797_ egd_top.BitStream_buffer.pc_reg\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4748_ _0731_ _0976_ _0347_ _0977_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4679_ _0587_ _0831_ _0832_ _2822_ _1391_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6418_ net160 _0251_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[6] sky130_fd_sc_hd__buf_12
X_6349_ net91 _0182_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[81\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3981_ _3069_ _2791_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__2724_ clknet_0__2724_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2724_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5720_ _2357_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ net4 _0395_ _2317_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__mux2_1
X_5582_ _2284_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__clkbuf_1
X_4602_ _1171_ _3093_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4533_ _2874_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4464_ _0874_ _0742_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__nand2_1
X_4395_ _3133_ _0976_ _0575_ _0977_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3415_ _2832_ _2875_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__nor2_4
X_6134_ _2565_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__inv_2
X_3346_ _2883_ _2764_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__nor2_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _2634_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__inv_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _1403_ _0811_ _1725_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3277_ _2827_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__clkbuf_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6225__91 clknet_1_1__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
X_5918_ _2491_ _2481_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _2431_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3200_ _2768_ egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\] vssd1
+ vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__and3_2
X_4180_ _2965_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3964_ _3024_ _2806_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5703_ net10 _0389_ _2334_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__mux2_1
X_3895_ _0430_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _0614_
+ sky130_fd_sc_hd__nand2_1
X_5634_ _2311_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ _0967_ _2881_ _0968_ _2943_ _2270_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__a221oi_1
X_4516_ _1224_ _1226_ _1228_ _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__and4_1
X_5496_ _0349_ _2911_ _3144_ _2916_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__o22ai_1
X_4447_ _0844_ _2987_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__nand2_1
X_4378_ _0933_ _0583_ _0934_ _0871_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__a22o_1
X_6117_ _2684_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__inv_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _2877_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__buf_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _2565_ _2589_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6204__72 clknet_1_1__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
XFILLER_0_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3680_ _0390_ _0393_ _0396_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5350_ _0797_ _2820_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__nand2_1
X_6274__136 clknet_1_0__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
X_4301_ _3058_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__clkinv_4
X_5281_ _0883_ _0412_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__nand2_1
X_4232_ _0384_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__clkbuf_4
X_4163_ _0871_ _0872_ _0657_ _0873_ _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__a221oi_1
X_4094_ _2982_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4996_ _1668_ _1677_ _1691_ _1706_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__and4_1
X_3947_ _2976_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _0665_
+ sky130_fd_sc_hd__nand2_1
X_3878_ _0394_ _2935_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__nand2_1
X_5617_ net4 _3010_ _2299_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5548_ _0925_ _0638_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__nand2_1
X_5479_ _0816_ _2806_ _0817_ _2874_ _2184_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__a221oi_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout50 net51 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_4
XFILLER_0_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4850_ _0974_ egd_top.BitStream_buffer.BS_buffer\[46\] _0975_ _2931_ _1561_ vssd1
+ vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3801_ _3020_ _2810_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__nand2_1
X_4781_ _1491_ _1492_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3732_ _0416_ _0426_ _0437_ _0451_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__and4_1
X_3663_ _0382_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0383_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6451_ net193 _0284_ net38 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6382_ net124 _0215_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[74\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5402_ _1171_ _0404_ _0480_ _0408_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5333_ _0463_ _0961_ _0962_ _2830_ _2040_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__a221oi_1
X_3594_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5264_ _1017_ _2854_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4215_ _0371_ _0930_ _0931_ _0553_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__a22o_1
X_5195_ _0859_ _0405_ _3091_ _0409_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__o22ai_1
X_4146_ _2929_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__clkbuf_8
X_4077_ _3058_ _0787_ _0402_ _0788_ _0793_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4979_ _1688_ _1689_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6195__63 clknet_1_0__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__inv_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6305__165 clknet_1_1__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__inv_2
XFILLER_0_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4000_ _0717_ _3131_ _0575_ _3135_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__o22ai_1
X_5951_ _2523_ _2527_ _2509_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _2804_ _0810_ _3066_ _0809_ _1612_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ _2458_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__inv_2
X_4833_ _0653_ _3110_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4764_ _1465_ _1469_ _1473_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6326__16 clknet_1_1__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__inv_2
X_3715_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6434_ net176 _0267_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_4695_ _0867_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _1408_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3646_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ net107 _0198_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3577_ _3125_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__buf_4
X_5316_ egd_top.BitStream_buffer.BS_buffer\[78\] _0930_ _0931_ _0657_ vssd1 vssd1
+ vccd1 vccd1 _2024_ sky130_fd_sc_hd__a22o_1
X_6296_ clknet_1_0__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__buf_1
X_5247_ _0820_ _2828_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__nand2_1
X_5178_ _3100_ _3040_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__nand2_1
X_4129_ _0546_ _0843_ _0845_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6159__30 clknet_1_1__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__inv_2
XFILLER_0_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6174__44 clknet_1_0__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__inv_2
X_3500_ _2845_ _2961_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__nand2_1
X_4480_ _0341_ _3126_ _0343_ _3123_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__a221oi_1
X_3431_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _2565_ _2708_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__nor2_1
X_3362_ _2884_ _2910_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__nand2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _1000_ _0945_ _0946_ _2931_ _1810_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__a221oi_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _2648_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__inv_2
X_3293_ egd_top.BitStream_buffer.pc\[0\] _2841_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__nand2_4
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _2867_ _0395_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5934_ _2498_ _2503_ _2510_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__nand3_2
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5865_ _2440_ _2441_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__nand2_1
X_4816_ _0877_ _2939_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__nand2_1
X_5796_ egd_top.BitStream_buffer.pc_reg\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__or2_1
X_4747_ _0967_ _2874_ _0968_ _0469_ _1459_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4678_ _1389_ _1390_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3629_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
X_6417_ net159 _0250_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_6348_ net90 _0181_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[82\]
+ sky130_fd_sc_hd__dfrtp_4
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[7] sky130_fd_sc_hd__buf_12
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__inv_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2723_ clknet_0__2723_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2723_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5650_ _2320_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
X_4601_ _3100_ _2887_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__nand2_1
X_5581_ net5 _0777_ _2281_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__mux2_1
X_4532_ _1193_ _0903_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__nand3_1
X_4463_ egd_top.BitStream_buffer.BS_buffer\[54\] _0863_ _0864_ _3119_ _1177_ vssd1
+ vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3414_ _2962_ _2816_ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__nand2_1
X_4394_ _0967_ _0777_ _0968_ _1011_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6133_ _2700_ _2554_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__nand2_1
X_3345_ _2893_ _2872_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__nand2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6064_ _2632_ _2633_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__nand2_1
X_3276_ net8 _2826_ _2797_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__mux2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _0812_ _2913_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__nand2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5917_ _2493_ _2466_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5848_ net12 _0583_ _2420_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5779_ _2389_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3963_ _3022_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _0681_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5702_ _2347_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
X_3894_ _0428_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _0613_
+ sky130_fd_sc_hd__nand2_1
X_5633_ net11 _2922_ _2299_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5564_ _0888_ _0969_ _1075_ _0971_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__o22ai_1
X_4515_ _0974_ _0336_ _0975_ _3146_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5495_ _0742_ _2839_ _2846_ _0871_ _2200_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__a221oi_1
X_4446_ _1150_ _1154_ _1156_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__and4_1
X_6251__115 clknet_1_0__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
X_4377_ _0656_ _0930_ _0931_ _0709_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__a22o_1
X_6116_ _2447_ _2516_ _2451_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__o21ai_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _2876_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__and3_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _2815_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__clkbuf_1
X_6047_ _2621_ _2554_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4300_ _0625_ _0781_ _3053_ _0782_ _1015_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__a221oi_1
X_5280_ _0892_ _0495_ _0893_ _0871_ _1987_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ _0947_ _0389_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nand2_1
X_4162_ _0876_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__nand2_1
X_4093_ _2989_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__clkbuf_4
X_4995_ _1694_ _1698_ _1702_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__and4_2
X_3946_ _2973_ _3143_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3877_ _0391_ _3142_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5616_ _2302_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__clkbuf_1
X_5547_ _3034_ _0933_ _3048_ _0934_ _2252_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__a221oi_1
X_5478_ _2182_ _2183_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__nand2_1
X_4429_ _0804_ _2824_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__nand2_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout40 net41 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_4
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout51 net52 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_2
XFILLER_0_91_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4780_ _0804_ _0458_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__nand2_1
X_3800_ _0517_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__nor2_1
X_3731_ _0442_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ _2864_ _2937_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__and2_1
X_6450_ net192 _0283_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3593_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__clkbuf_8
X_6381_ net123 _0214_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[75\]
+ sky130_fd_sc_hd__dfrtp_4
X_5401_ _2064_ _2078_ _2090_ _2107_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__and4_1
X_5332_ _0543_ _0963_ _3129_ _0964_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__o22ai_1
X_5263_ _2858_ _0920_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5194_ _1896_ _1898_ _1900_ _1902_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__and4_1
X_4214_ _0370_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4145_ _0847_ _0853_ _0856_ _0861_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ _0789_ _0790_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4978_ _1017_ _0446_ _1126_ _0449_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3929_ _2938_ _0346_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _2526_ _2508_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__nand2_1
X_4901_ _1287_ _0811_ _1611_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5881_ _2456_ _2457_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__nand2_1
X_4832_ _3118_ _0389_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4763_ _1474_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6502_ net76 _0328_ net39 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dfrtp_2
X_3714_ _2895_ _2837_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__and2_1
X_4694_ _0865_ _0336_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__nand2_1
X_6433_ net175 _0266_ net41 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3645_ _0358_ _0360_ _0362_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__and4_1
X_6364_ net106 _0197_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_3576_ _2927_ _2909_ vssd1 vssd1 vccd1 vccd1 _3125_ sky130_fd_sc_hd__and2_1
X_5315_ _2008_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__and2_1
X_5246_ _0818_ _0777_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5177_ _0392_ _0907_ _0371_ _0908_ _1885_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__a221oi_1
X_4128_ _0844_ _0610_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__nand2_1
X_4059_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3430_ _2942_ _2955_ _2968_ _2978_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__and4_1
X_3361_ _2909_ vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__clkbuf_4
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080_ _2639_ _2644_ _2615_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__a21oi_2
X_5100_ _1808_ _1809_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__nand2_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3292_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__inv_2
X_5031_ _2943_ _0840_ _2887_ _0842_ _1740_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__a221oi_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _2508_ _2509_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__nand2_1
X_5864_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1 vccd1
+ _2441_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4815_ _0874_ _0420_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__nand2_1
X_5795_ _2398_ _2399_ _2400_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__a21bo_2
X_4746_ _0561_ _0969_ _3075_ _0971_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4677_ _0835_ _0625_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3628_ _2946_ _2937_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__nand2_1
X_6416_ net158 _0249_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6347_ net89 _0180_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[83\]
+ sky130_fd_sc_hd__dfrtp_4
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 la_data_out_18_16[0] sky130_fd_sc_hd__buf_12
X_3559_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__inv_2
X_5229_ _1936_ _1937_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2722_ clknet_0__2722_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2722_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4600_ egd_top.BitStream_buffer.BS_buffer\[57\] _0907_ _3139_ _0908_ _1313_ vssd1
+ vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__a221oi_2
X_5580_ _2283_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4531_ _1206_ _1222_ _1231_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__and4_1
X_4462_ _1175_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__nand2_1
X_3413_ _2864_ _2961_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__and2_1
X_4393_ _0543_ _0969_ _0347_ _0971_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6132_ _2695_ _2699_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__nand2_1
X_3344_ _2892_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__buf_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _2505_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1
+ vccd1 _2633_ sky130_fd_sc_hd__nand2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5014_ _1713_ _1716_ _1719_ _1723_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__and4_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5916_ _2492_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5847_ _2430_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
X_5778_ net11 _3058_ _2377_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4729_ _0638_ _0922_ _0583_ _0921_ _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3962_ _3020_ _2812_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5701_ net11 _0385_ _2335_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3893_ _0606_ _0608_ _0609_ _0611_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__and4_1
X_5632_ _2310_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
X_5563_ _0464_ _0961_ _0962_ _2848_ _2268_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__a221oi_1
X_4514_ _0349_ _0976_ _0731_ _0977_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5494_ _3154_ _2853_ _2199_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__o21ai_1
X_4445_ _0920_ _0831_ _0832_ _2818_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__a221oi_2
X_4376_ _0875_ _0921_ _0607_ _0922_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__a221oi_1
X_6115_ _2595_ _2663_ _2682_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__nand3_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _2875_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__inv_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ net14 _2814_ _2798_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__mux2_1
X_6046_ _2617_ _2620_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__nand2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ net18 vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4230_ _0382_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__clkbuf_4
X_4161_ _0877_ _0336_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ _2986_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__clkbuf_4
X_4994_ _1703_ _1704_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3945_ _2971_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _0663_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5615_ net5 _2993_ _2299_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__mux2_1
X_3876_ _0388_ _2951_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6210__77 clknet_1_1__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
X_5546_ _0495_ _0930_ _0931_ _1000_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__a22o_1
X_5477_ _0820_ _0625_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4428_ _0802_ _2791_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__nand2_1
X_4359_ _0389_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__inv_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _2600_ _2603_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout52 net19 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_4
Xfanout41 net42 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6280__142 clknet_1_0__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3730_ _0444_ _0446_ _0447_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3661_ _0380_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _0381_
+ sky130_fd_sc_hd__nand2_1
X_6380_ net122 _0213_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[76\]
+ sky130_fd_sc_hd__dfrtp_4
X_3592_ _3140_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__clkbuf_2
X_5400_ _2094_ _2098_ _2102_ _2106_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__and4_1
X_5331_ _2822_ _0954_ _2820_ _0955_ _2038_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5262_ _0402_ _0848_ _2913_ _0849_ _1969_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5193_ _0974_ _2926_ _0975_ _0346_ _1901_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__a221oi_1
X_4213_ _0368_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__clkbuf_4
X_4144_ _2980_ _0857_ _3097_ _0858_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _0791_ _3030_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4977_ _0439_ _2987_ _0441_ _3034_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3928_ _2934_ _0341_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nand2_1
X_3859_ _0576_ _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5529_ _2233_ _2234_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4900_ _0812_ _2922_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nand2_1
X_5880_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] vssd1 vssd1 vccd1 vccd1
+ _2457_ sky130_fd_sc_hd__inv_2
X_4831_ _0333_ _3126_ _3143_ _3123_ _1542_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4762_ _0686_ _0446_ _0772_ _0449_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6501_ net75 _0327_ net39 vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dfrtp_2
X_3713_ _0432_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _0433_
+ sky130_fd_sc_hd__nand2_1
X_4693_ _1396_ _1399_ _1402_ _1405_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__and4_1
X_6432_ net174 _0265_ net41 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_3644_ _0363_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _0364_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3575_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__clkbuf_8
X_6363_ net105 _0196_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5314_ _2011_ _2014_ _2018_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__and4_1
X_5245_ _2810_ _0810_ _0330_ _0809_ _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5176_ _1185_ _3110_ _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__o21ai_1
X_6287__148 clknet_1_0__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__inv_2
X_4127_ _2903_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__clkbuf_4
X_4058_ _0720_ _0735_ _0755_ _0775_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6331__21 clknet_1_0__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__inv_2
X_3360_ _2768_ _2834_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2909_
+ sky130_fd_sc_hd__and3_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3291_ _2839_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__buf_4
X_5030_ _3008_ _0843_ _1739_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__o21ai_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5932_ _2488_ _2481_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5863_ _2438_ _2439_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5794_ egd_top.BitStream_buffer.pc_reg\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ egd_top.BitStream_buffer.BS_buffer\[57\] _0863_ _0864_ egd_top.BitStream_buffer.BS_buffer\[55\]
+ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__a221oi_2
X_4745_ _3105_ _0961_ _0962_ _0656_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4676_ _0833_ _2816_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3627_ _0346_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
X_6415_ net157 _0248_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_3558_ _3091_ _3093_ _3098_ _3102_ _3106_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__o2111a_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 la_data_out_18_16[1] sky130_fd_sc_hd__buf_12
X_6346_ net88 _0179_ net51 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[84\]
+ sky130_fd_sc_hd__dfrtp_4
X_6180__49 clknet_1_1__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__inv_2
X_3489_ _3036_ _3037_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__nand2_1
X_5228_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1
+ vccd1 _1937_ sky130_fd_sc_hd__nand2_1
X_5159_ _0874_ _0477_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2721_ clknet_0__2721_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2721_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4530_ _1233_ _1237_ _1241_ _1244_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4461_ _0867_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _1176_
+ sky130_fd_sc_hd__nand2_1
X_3412_ _2960_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__buf_2
X_4392_ _2957_ _0961_ _0962_ _0435_ _1107_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6131_ _2696_ _2698_ _2514_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3343_ _2765_ egd_top.BitStream_buffer.pc\[2\] _2868_ vssd1 vssd1 vccd1 vccd1 _2892_
+ sky130_fd_sc_hd__and3_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _2481_ _2499_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] vssd1
+ vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__o21ai_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _2825_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5013_ _2804_ _0800_ _0801_ _2826_ _1722_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__a221oi_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5915_ _2491_ _2476_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5846_ net13 _0742_ _2420_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777_ _2388_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4728_ _1439_ _1440_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4659_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6216__83 clknet_1_0__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
XFILLER_0_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _0677_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5700_ _2346_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3892_ _0424_ _0610_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5631_ net12 _2920_ _2299_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5562_ _3129_ _0963_ _0717_ _0964_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__o22ai_1
X_4513_ _0967_ _1011_ _0968_ _0886_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a221oi_1
X_5493_ _2857_ _0587_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__nand2_1
X_4444_ _1157_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__nand2_1
X_4375_ _1089_ _1090_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__nand2_1
X_6114_ _2634_ _2667_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__nor2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _2763_ _2841_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__nand2_4
X_6045_ _2593_ _2590_ _2619_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__nand3_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__buf_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ net17 vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5829_ _2421_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4160_ _2973_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4091_ _0786_ _0794_ _0799_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _0933_ _0477_ _0934_ _0638_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__a22o_1
X_3944_ _2969_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0662_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3875_ _0590_ _0591_ _0592_ _0593_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5614_ _2301_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5545_ _2236_ _2250_ vssd1 vssd1 vccd1 vccd1 _2251_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ _0818_ _0886_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4427_ _1140_ _3065_ _3064_ _0796_ _1141_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _1028_ _1042_ _1055_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__and4_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _1005_ _0446_ _0465_ _0449_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o22ai_1
X_3309_ _2857_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__clkbuf_4
X_6028_ _2601_ _2602_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__nand2_1
Xfanout42 net46 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_2
XFILLER_0_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3660_ _2864_ _2837_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__and2_1
X_3591_ _2884_ _2836_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__and2_1
X_5330_ _3154_ _0956_ _1488_ _0958_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5261_ _3008_ _0850_ _1968_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__o21ai_1
X_4212_ _0920_ _0921_ _0420_ _0922_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__a221oi_1
X_5192_ _0730_ _0976_ _0543_ _0977_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ _0859_ _2912_ _3091_ _2917_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__o22ai_1
X_4074_ _3033_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4976_ _0463_ _0996_ _2959_ _0997_ _1686_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__a221oi_1
X_3927_ _0632_ _0635_ _0640_ _0644_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3858_ _0352_ egd_top.BitStream_buffer.BS_buffer\[127\] _0353_ egd_top.BitStream_buffer.BS_buffer\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3789_ _2989_ _3058_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__nand2_1
X_5528_ _0957_ _0445_ _1017_ _0448_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__o22ai_1
X_5459_ _2164_ _2165_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__nand2_1
X_6264__127 clknet_1_1__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
X_6186__55 clknet_1_1__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__inv_2
XFILLER_0_52_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4830_ _0888_ _3131_ _3075_ _3135_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__o22ai_1
X_4761_ _0439_ _0610_ _0441_ _0443_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__a22o_1
X_6500_ net74 _0326_ net39 vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfrtp_4
X_3712_ _2884_ _2851_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4692_ _3127_ _0857_ _3124_ _0858_ _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6431_ net173 _0264_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_3643_ _2864_ _2852_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6362_ net104 _0195_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_5313_ _2019_ _2020_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__nor2_1
X_3574_ _3122_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__buf_4
X_5244_ _0334_ _0811_ _1951_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5175_ _3118_ _3142_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__nand2_1
X_4126_ _2894_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4057_ _0760_ _0765_ _0770_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4959_ _2816_ _0954_ _2814_ _0955_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _2838_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6247__111 clknet_1_1__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_0_18_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5931_ _2504_ _2507_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5862_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1 vccd1
+ _2439_ sky130_fd_sc_hd__inv_2
X_5793_ egd_top.BitStream_buffer.pc_reg\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__or2_1
X_4813_ _1523_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__nand2_1
X_4744_ _0970_ _0963_ _0574_ _0964_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4675_ _0824_ _2980_ _0825_ _3097_ _1387_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__a221oi_1
X_6165__36 clknet_1_1__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__inv_2
X_3626_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__buf_4
X_6414_ net156 _0247_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3557_ _3104_ _3105_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__nand2_1
X_6345_ net87 _0178_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[85\]
+ sky130_fd_sc_hd__dfrtp_4
X_3488_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__clkbuf_8
X_5227_ _1934_ _1935_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__nand2_1
X_5158_ _0389_ _0863_ _0864_ _3115_ _1866_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__a221oi_1
X_4109_ _3009_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__clkbuf_4
X_5089_ _1797_ _1798_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__nand2_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2720_ clknet_0__2720_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2720_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _0865_ _0333_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_1
X_4391_ _0349_ _0963_ _0731_ _0964_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__o22ai_1
X_3411_ egd_top.BitStream_buffer.pc\[6\] egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6130_ _2648_ _2697_ _2690_ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__o21ai_1
X_3342_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__inv_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _2603_ _2569_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__nand2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ net9 _2824_ _2797_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__mux2_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _1720_ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__nand2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5914_ _2488_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__inv_6
XFILLER_0_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5845_ _2429_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5776_ net12 _2990_ _2377_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__mux2_1
X_4727_ _0925_ _0742_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4658_ _0330_ _0787_ _2913_ _0788_ _1370_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__a221oi_1
X_3609_ _2767_ _2985_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4589_ _3011_ _0882_ _1299_ _1300_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_12_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ _3014_ _0402_ _3016_ _2863_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__a22o_1
X_3891_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _2309_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
X_5561_ _2826_ _0954_ _2824_ _0955_ _2266_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4512_ _3108_ _0969_ _0574_ _0971_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__o22ai_1
X_5492_ _2920_ _0848_ _3097_ _0849_ _2197_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4443_ _0835_ _2828_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__nand2_1
X_4374_ _0925_ _0920_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__nand2_1
X_6113_ _2509_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__inv_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__clkbuf_8
X_3256_ _2813_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__clkbuf_1
X_6044_ _2618_ _2512_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__nand2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _2754_ _2755_ _2756_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5828_ net7 _0495_ _2420_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5759_ _2379_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4090_ _3066_ _0800_ _0801_ _2812_ _0806_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__a221oi_1
X_4992_ egd_top.BitStream_buffer.BS_buffer\[75\] _0930_ _0931_ egd_top.BitStream_buffer.BS_buffer\[78\]
+ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _2956_ _0656_ _2958_ _0657_ _0660_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a221oi_1
X_3874_ _0384_ _0389_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5613_ net6 _3007_ _2299_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6312__3 clknet_1_1__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__inv_2
X_5544_ _2239_ _2242_ _2246_ _2249_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__and4_1
X_5475_ _2800_ _0809_ _2814_ _0810_ _2180_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4426_ _0797_ _2804_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__nand2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _1059_ _1063_ _1068_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__and4_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__inv_2
X_3308_ _2856_ _2837_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__and2_1
X_3239_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__buf_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _2505_ _2441_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout43 net44 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_4
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6241__106 clknet_1_1__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3590_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5260_ _2867_ _0378_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__nand2_1
X_4211_ _0924_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nand2_1
X_5191_ _0967_ _0841_ _0968_ _3101_ _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__a221oi_1
X_4142_ _0395_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__inv_2
X_4073_ _3032_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4975_ _1684_ _1685_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _0642_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__nor2_1
X_3857_ _0574_ _0348_ _0575_ _0350_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3788_ _2986_ _3034_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nand2_1
X_5527_ _0438_ _3037_ _0440_ _3053_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__a22o_1
X_5458_ net221 egd_top.BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1
+ vccd1 _2165_ sky130_fd_sc_hd__nand2_1
X_4409_ _0439_ _2904_ _0441_ _0477_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__a22o_1
X_5389_ _0877_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _2096_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4760_ _2859_ _0996_ _2848_ _0997_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__a221oi_1
X_3711_ _0430_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _0431_
+ sky130_fd_sc_hd__nand2_1
X_4691_ _1403_ _2912_ _0859_ _2917_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__o22ai_1
X_6430_ net172 _0263_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_3642_ _0361_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _0362_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6361_ net103 _0194_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3573_ _2946_ _2909_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__and2_1
X_5312_ _1417_ _3130_ _0561_ _3134_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5243_ _0812_ _3097_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__nand2_1
X_5174_ _3146_ _3126_ _3132_ _3123_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__a221oi_1
X_4125_ _2900_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__clkbuf_4
X_4056_ _0771_ _0773_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4958_ _0789_ _0956_ _1140_ _0958_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_46_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4889_ _0791_ _3153_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3909_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] vssd1 vssd1
+ vccd1 vccd1 _0628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5930_ _2505_ _2506_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5861_ _2437_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1
+ vccd1 _2438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5792_ _2762_ _2397_ _2396_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__o21ai_4
X_4812_ _0867_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _1524_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4743_ _2812_ _0954_ _2810_ _0955_ _1455_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4674_ _0403_ _0826_ _0756_ _0827_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__o22ai_1
X_6413_ net155 _0246_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_3625_ _0339_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__nor2_1
X_3556_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__clkbuf_8
X_6344_ net86 _0177_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[86\]
+ sky130_fd_sc_hd__dfrtp_4
X_6293__154 clknet_1_1__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__inv_2
X_5226_ _0551_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3487_ _2964_ _2985_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__and2_1
X_5157_ _1864_ _1865_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__nand2_1
X_4108_ _3016_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__clkbuf_4
X_5088_ _0999_ _0583_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__nand2_1
X_4039_ _3015_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4390_ _2806_ _0954_ _2804_ _0955_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__a221oi_2
X_3410_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__clkbuf_8
X_6170__40 clknet_1_1__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__inv_2
X_3341_ _2863_ _2867_ _2873_ _2874_ _2889_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _2622_ _2623_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__nand2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__clkbuf_8
X_5011_ _0804_ _0777_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__nand2_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5913_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] _2489_ vssd1 vssd1 vccd1
+ vccd1 _2490_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5844_ net14 _0587_ _2420_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5775_ _2387_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4726_ _0923_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _1439_
+ sky130_fd_sc_hd__or2b_1
X_6301__161 clknet_1_0__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__inv_2
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4657_ _0567_ _0790_ _1369_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__o21ai_1
X_3608_ _2884_ _2996_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4588_ _1301_ _0889_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__or2_1
X_3539_ _3087_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _3088_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5209_ _0925_ _0607_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6207__74 clknet_1_0__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
X_3890_ _0422_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0609_
+ sky130_fd_sc_hd__nand2_1
X_6222__88 clknet_1_0__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
X_5560_ _0723_ _0956_ _1717_ _0958_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__o22ai_2
X_4511_ _0371_ _0961_ _0962_ _2957_ _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__a221oi_1
X_5491_ _3011_ _0850_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4442_ _0833_ _2812_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ _0923_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _1089_
+ sky130_fd_sc_hd__or2b_1
X_6112_ _2656_ _2675_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _2870_ _2872_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__and2_1
X_3255_ net15 _2812_ _2798_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__mux2_1
X_6043_ _2605_ _2614_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__nand2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ egd_top.BitStream_buffer.pc_previous\[5\] egd_top.BitStream_buffer.pc_previous\[4\]
+ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5827_ _2419_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__buf_4
XFILLER_0_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5758_ net6 _0610_ _2377_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__mux2_1
X_4709_ _1420_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nand2_1
X_5689_ net2 egd_top.BitStream_buffer.BS_buffer\[53\] _2335_ vssd1 vssd1 vccd1 vccd1
+ _2341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4991_ _0937_ _0371_ _3105_ _0938_ _1701_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__a221oi_1
X_3942_ _0658_ _0659_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3873_ _0382_ _3115_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5612_ _2300_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5543_ _2247_ _2248_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5474_ _0337_ _0811_ _2179_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4425_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__inv_2
X_4356_ _0892_ _0553_ _0893_ _1000_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__a221oi_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _2832_ _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__nor2_4
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _0439_ _0607_ _0441_ _2904_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__a22o_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _2516_ _2445_ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__nand2_1
X_3238_ _2801_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_1
X_3169_ _2733_ _2736_ net32 _2740_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout44 net45 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_4
X_6201__69 clknet_1_1__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__inv_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4210_ _0925_ _0926_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5190_ _2952_ _0969_ _0561_ _0971_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__o22ai_1
X_4141_ _2921_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__buf_4
X_4072_ _2990_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4974_ _0999_ _0742_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3925_ _2919_ _2913_ _2921_ _2980_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3856_ _2931_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3787_ _3097_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__inv_2
X_5526_ egd_top.BitStream_buffer.BS_buffer\[81\] _0996_ _0830_ _0997_ _2231_ vssd1
+ vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__a221oi_1
X_5457_ _2162_ _2163_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__nand2_1
X_4408_ _3105_ _0996_ _2859_ _0997_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__a221oi_1
X_5388_ _0874_ _0610_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4339_ _1045_ _1048_ _1051_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6009_ _2456_ _2584_ _2494_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3710_ _2899_ _2837_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4690_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _2895_ _2852_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3572_ _3108_ _3110_ _3113_ _3116_ _3120_ vssd1 vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__o2111a_1
X_6360_ net102 _0193_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_5311_ _3122_ egd_top.BitStream_buffer.BS_buffer\[46\] _3125_ _3132_ vssd1 vssd1
+ vccd1 vccd1 _2019_ sky130_fd_sc_hd__a22o_1
X_5242_ _1939_ _1942_ _1945_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__and4_2
X_5173_ _1301_ _3131_ _3129_ _3135_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__o22ai_1
X_4124_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__clkbuf_8
Xinput1 la_data_in_47_32[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4055_ _0772_ _0446_ _2849_ _0449_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4957_ _1657_ _1660_ _1663_ _1667_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__and4_1
X_3908_ _0542_ _0624_ _0457_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__a31o_1
X_4888_ _0469_ _0781_ _3070_ _0782_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__a221oi_2
X_3839_ _3118_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _0558_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6191__60 clknet_1_0__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__inv_2
X_6489_ net63 _0322_ net36 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dfrtp_4
X_5509_ _2213_ _2214_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2719_ clknet_0__2719_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2719_
+ sky130_fd_sc_hd__clkbuf_16
X_5860_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1 vccd1
+ _2437_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _0865_ _3146_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5791_ _2395_ _2396_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__nand2_2
X_4742_ _0526_ _0956_ _0795_ _0958_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4673_ _0816_ _3153_ _0817_ _2826_ _1385_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3624_ _0340_ _0341_ _0342_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__a22o_1
X_6412_ net154 _0245_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6343_ net85 _0176_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[87\]
+ sky130_fd_sc_hd__dfrtp_2
X_3555_ _3103_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__buf_4
X_3486_ _3033_ _3034_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__nand2_1
X_5225_ _1881_ _0903_ _1933_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5156_ _0867_ _0385_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__nand2_1
X_4107_ _3014_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__clkbuf_4
X_5087_ _0428_ _0920_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__nand2_1
X_4038_ _2920_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6228__94 clknet_1_1__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _2558_ net18 _2559_ _2758_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__a31o_2
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6156__27 clknet_1_0__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__inv_2
XFILLER_0_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6277__139 clknet_1_1__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3340_ _2882_ _2888_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__nand2_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _0802_ _2808_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__nand2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _2823_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__clkbuf_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5912_ _2466_ _2482_ _2488_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5843_ _2428_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5774_ net13 _3053_ _2377_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4725_ _1427_ _1430_ _1433_ _1437_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__and4_1
X_4656_ _0791_ _3058_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__nand2_1
X_3607_ _3151_ _3152_ _3154_ _3155_ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__o22ai_1
X_4587_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__inv_2
X_3538_ _3086_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__clkbuf_4
X_3469_ _3014_ _3015_ _3016_ _3017_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6257_ clknet_1_0__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__buf_1
X_5208_ _1905_ _1909_ _1913_ _1916_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__and4_1
X_5139_ _0835_ _2874_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4510_ _0575_ _0963_ _0970_ _0964_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5490_ _2866_ _0343_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4441_ _0824_ _2922_ _0825_ _2913_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__a221oi_1
X_6111_ _2646_ _2565_ _2679_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__o21ai_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _1077_ _1080_ _1083_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__and4_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _2871_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__clkbuf_4
X_3254_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__buf_4
X_6042_ _2594_ _2616_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__nand2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ egd_top.BitStream_buffer.pc_previous\[3\] egd_top.BitStream_buffer.pc_previous\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5826_ _2773_ egd_top.BitStream_buffer.buffer_index\[5\] _2775_ _2793_ vssd1 vssd1
+ vccd1 vccd1 _2419_ sky130_fd_sc_hd__or4b_4
XFILLER_0_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5757_ _2378_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4708_ _0897_ _2959_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__nand2_1
X_5688_ _2340_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
X_4639_ _0412_ _0987_ _3101_ _0989_ _1352_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6309_ clknet_1_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__buf_1
XFILLER_0_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6308__168 clknet_1_1__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__inv_2
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4990_ _1699_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3941_ _2965_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _0659_
+ sky130_fd_sc_hd__nand2_1
X_3872_ _0380_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _0591_
+ sky130_fd_sc_hd__nand2_1
X_5611_ net7 _2887_ _2299_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__mux2_1
X_5542_ _1647_ _3130_ _0904_ _3134_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5473_ _0812_ _2907_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__nand2_1
X_4424_ _3153_ _0787_ _2920_ _0788_ _1138_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4355_ _1069_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__nand2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _2763_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__nand2_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _0656_ _0996_ _0709_ _0997_ _1002_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__a221oi_1
X_3237_ net6 _2800_ _2798_ vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__mux2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _2508_ _2522_ _2569_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__nand3_1
X_3168_ _2739_ _2736_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6198__66 clknet_1_0__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__inv_2
Xfanout45 net46 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_4
X_5809_ _2410_ _2405_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _2919_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__buf_4
X_4071_ _3039_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__buf_4
X_4973_ _0428_ _0926_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3924_ _0641_ _2912_ _0506_ _2917_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6329__19 clknet_1_1__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__inv_2
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3855_ _3112_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__inv_2
X_3786_ _0488_ _0494_ _0499_ _0504_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__and4_1
X_5525_ _2229_ _2230_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ _2943_ _0456_ _2790_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__o21a_1
X_4407_ _1121_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_1
X_5387_ _0392_ _0863_ _0864_ _0389_ _2093_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__a221oi_2
X_4338_ _3097_ _0857_ _3090_ _0858_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ _0981_ _3007_ _0982_ _2993_ _0985_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__a221oi_1
X_6008_ _2455_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1
+ vccd1 vccd1 _2584_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6177__47 clknet_1_0__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__inv_2
XFILLER_0_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _0359_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0360_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3571_ _3118_ _3119_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__nand2_1
X_5310_ _1066_ _3076_ _2015_ _2016_ _2017_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5241_ _2808_ _0800_ _0801_ _0458_ _1948_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__a221oi_1
X_5172_ _1837_ _1851_ _1863_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__and4_1
X_4123_ _2896_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__clkbuf_4
Xinput2 la_data_in_47_32[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_4
X_4054_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _0492_ _3077_ _1664_ _1665_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__o2111a_1
X_3907_ _0625_ _0456_ _2789_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__o21ai_1
X_4887_ egd_top.BitStream_buffer.BS_buffer\[4\] _0783_ _0784_ _2874_ vssd1 vssd1 vccd1
+ vccd1 _1598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3838_ _3114_ _0385_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5508_ _0897_ _0920_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__nand2_1
X_3769_ _0346_ _2929_ _2930_ _2939_ _0487_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__a221oi_2
X_6488_ net62 _0321_ net38 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_valid_n
+ sky130_fd_sc_hd__dfstp_1
X_5439_ _0937_ _0709_ _2830_ _0938_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__a221oi_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2718_ clknet_0__2718_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2718_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4810_ _1512_ _1515_ _1518_ _1521_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5790_ egd_top.BitStream_buffer.pc_reg\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4741_ _1442_ _1445_ _1449_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__and4_1
X_4672_ _1383_ _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6411_ net153 _0244_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_3623_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6254__118 clknet_1_0__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
X_6342_ net84 _0175_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[88\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3554_ _2893_ _2837_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__and2_2
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3485_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__buf_4
X_5224_ _1894_ _1903_ _1917_ _1932_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5155_ _0865_ _2931_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__nand2_1
X_4106_ _0816_ _3053_ _0817_ _2818_ _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__a221oi_1
X_5086_ _2993_ _0987_ _0412_ _0989_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__a221oi_1
X_4037_ _0740_ _0744_ _0749_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ net17 _2759_ _2514_ _2564_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__a31o_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4939_ _0895_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _1650_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_40 _3101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ net10 _2822_ _2797_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__mux2_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5911_ _2485_ _2487_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__nand2_4
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5842_ net15 _0875_ _2420_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5773_ _2386_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ _1075_ _3077_ _1434_ _1435_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_31_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4655_ _0886_ _0781_ _3066_ _0782_ _1367_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3606_ _2845_ _2985_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4586_ _0885_ _0988_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__nand2_1
X_3537_ _2899_ _2937_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__and2_1
X_3468_ egd_top.BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__buf_4
X_5207_ _1914_ _1915_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__nor2_1
X_3399_ _2947_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _2948_
+ sky130_fd_sc_hd__nand2_1
X_5138_ _0833_ _2824_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__nand2_1
X_5069_ _3087_ _3139_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6237__102 clknet_1_0__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XFILLER_0_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4440_ _0757_ _0826_ _0403_ _0827_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_0_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6110_ _2676_ _2554_ _2678_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__nand3_1
X_4371_ _0561_ _3077_ _1084_ _1085_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__o2111a_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _2768_ _2834_ _2835_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__and3_2
X_3253_ _2811_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__clkbuf_1
X_6041_ _2605_ _2614_ _2615_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__a21oi_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.pc_previous\[0\]
+ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__nand2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5825_ _2418_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5756_ net7 _0638_ _2377_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5687_ net3 _3119_ _2335_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__mux2_1
X_4707_ _0895_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _1420_
+ sky130_fd_sc_hd__nand2_1
X_4638_ _1350_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ _2993_ _0848_ _3015_ _0849_ _1282_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__a221oi_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3940_ _2962_ _2820_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3871_ _0377_ _0341_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nand2_1
X_5610_ _2298_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5541_ _3122_ _2939_ _3125_ _2931_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5472_ _2167_ _2170_ _2173_ _2177_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__and4_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4423_ _3067_ _0790_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__o21ai_1
X_4354_ _0897_ _0463_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand2_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _2853_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__clkbuf_4
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _2595_ _2569_ _2598_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__nand3_1
X_4285_ _0998_ _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__nand2_1
X_3236_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__buf_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3167_ net31 vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout35 net36 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_4
Xfanout46 net19 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5808_ egd_top.BitStream_buffer.pc_reg\[4\] _2404_ vssd1 vssd1 vccd1 vccd1 _2410_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5739_ net9 _2848_ _2352_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _3036_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__clkbuf_4
X_6289__150 clknet_1_0__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__inv_2
XFILLER_0_25_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4972_ _3007_ _0987_ _2943_ _0989_ _1682_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__a221oi_1
X_3923_ _3124_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3854_ _0571_ _0572_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3785_ _0500_ _0501_ _0502_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__and4_1
X_5524_ _0999_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _2230_
+ sky130_fd_sc_hd__nand2_1
X_5455_ _2108_ _0903_ _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4406_ _0999_ _0830_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__nand2_1
X_5386_ _2091_ _2092_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4337_ _1052_ _2912_ _2908_ _2917_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o22ai_1
X_4268_ _0983_ _0405_ _0984_ _0409_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__o22ai_1
X_3219_ _2786_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__clkbuf_1
X_6007_ _2451_ _2543_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__nor2_1
X_4199_ _0544_ _3084_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3570_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__buf_4
XFILLER_0_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _1946_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5171_ _1867_ _1871_ _1875_ _1879_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__and4_1
X_4122_ _0815_ _0823_ _0829_ _0838_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__and4_1
X_4053_ _0439_ egd_top.BitStream_buffer.BS_buffer\[92\] _0441_ egd_top.BitStream_buffer.BS_buffer\[93\]
+ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__a22o_1
Xinput3 la_data_in_47_32[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_4
XFILLER_0_59_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4955_ _3087_ _3142_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__nand2_1
X_3906_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4886_ _1596_ _1597_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__nand2_1
X_3837_ _3111_ _3119_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__nand2_1
X_3768_ _0485_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__nand2_1
X_5507_ _0895_ _0988_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__nand2_1
X_3699_ _2878_ _2851_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__and2_1
X_6487_ net61 _0320_ net46 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_5438_ _2143_ _2144_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__nand2_1
X_5369_ _2074_ _2075_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6182__51 clknet_1_1__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__inv_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2717_ clknet_0__2717_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2717_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4740_ _0495_ _0945_ _0946_ _3146_ _1452_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4671_ _0820_ _2818_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3622_ _2893_ _2910_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__and2_1
X_6410_ net152 _0243_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[46\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6341_ net83 _0174_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[89\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3553_ _3100_ _3101_ vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3484_ _2933_ _2985_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5223_ _1920_ _1924_ _1928_ _1931_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__and4_1
X_5154_ _1854_ _1857_ _1860_ _1862_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__and4_1
X_4105_ _0819_ _0821_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__nand2_1
X_5085_ _1793_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__nand2_1
X_4036_ _0750_ _0751_ _0752_ _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _2553_ _2554_ _2555_ _2563_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__a31o_1
X_4938_ _0757_ _0882_ _1645_ _1646_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__o2111a_1
X_4869_ _0947_ _0398_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__nand2_1
XANTENNA_41 egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_30 _2864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6219__85 clknet_1_0__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6234__99 clknet_1_0__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
XFILLER_0_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ _2486_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6315__6 clknet_1_1__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__inv_2
X_5841_ _2427_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6260__123 clknet_1_1__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
X_5772_ net14 _3037_ _2377_ vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__mux2_1
X_4723_ _3087_ _2951_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4654_ egd_top.BitStream_buffer.BS_buffer\[2\] _0783_ _0784_ _1011_ vssd1 vssd1 vccd1
+ vccd1 _1367_ sky130_fd_sc_hd__a22o_1
X_3605_ _3153_ vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__inv_2
X_4585_ _0883_ _1116_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nand2_1
X_3536_ _3082_ _3084_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6161__32 clknet_1_1__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__inv_2
X_3467_ _2893_ _2915_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__and2_1
X_5206_ _3154_ _0446_ _0526_ _0449_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__o22ai_1
X_3398_ _2946_ _2872_ vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__and2_1
X_5137_ _0824_ _3127_ _0825_ _3124_ _1845_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__a221oi_1
X_5068_ _3011_ _3084_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__or2_1
X_4019_ _0359_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0737_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2719_ _2719_ vssd1 vssd1 vccd1 vccd1 clknet_0__2719_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4370_ _3087_ _3115_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3321_ _2869_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ net16 _2810_ _2798_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__mux2_1
X_6040_ _2760_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__inv_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ egd_top.BitStream_buffer.pc_previous\[6\] vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__inv_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5824_ egd_top.BitStream_buffer.pc\[0\] net38 vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ _2376_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5686_ _2339_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4706_ _0407_ _0882_ _1415_ _1416_ _1418_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__o2111a_1
X_4637_ _0992_ _3002_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4568_ _3078_ _0850_ _1281_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__o21ai_1
X_3519_ _2878_ _2985_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__nand2_1
X_4499_ _0939_ _2974_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__nand2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _0586_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5540_ _1301_ _3076_ _2243_ _2244_ _2245_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__o2111a_1
X_5471_ _2812_ _0800_ _0801_ _0777_ _2176_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ _0791_ _3053_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4353_ _0895_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _1069_
+ sky130_fd_sc_hd__nand2_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _0999_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__nand2_1
X_3304_ _2767_ _2852_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__nand2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ _2596_ _2597_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__nand2_1
X_3235_ _2799_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__clkbuf_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _2732_ _2737_ _2738_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout36 net46 vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_4
Xfanout47 net51 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_4
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3999_ _3115_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__inv_2
X_5807_ _2409_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5738_ _2366_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5669_ net10 _3146_ _2316_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4971_ _1680_ _1681_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3922_ _3082_ _2894_ _0636_ _0637_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3853_ _0340_ _0343_ _0342_ _2974_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3784_ _2976_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _0503_
+ sky130_fd_sc_hd__nand2_1
X_5523_ _0427_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _2229_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5454_ _2137_ _2151_ _2160_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__and3_1
X_4405_ _0428_ _0495_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nand2_1
X_5385_ _0867_ _2951_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4336_ _2935_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4267_ _3017_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__inv_2
X_4198_ _0489_ _3080_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__or2_1
X_3218_ _2785_ net29 _2783_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__mux2_1
X_6006_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _2542_ vssd1 vssd1 vccd1
+ vccd1 _2582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6319__10 clknet_1_0__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__inv_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6334__24 clknet_1_0__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__inv_2
X_5170_ _0403_ _0882_ _1876_ _1877_ _1878_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__o2111a_1
X_4121_ _0830_ _0831_ _0832_ _2814_ _0837_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__a221oi_1
X_4052_ _0766_ _0767_ _0768_ _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__and4_1
Xinput4 la_data_in_47_32[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_4
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4954_ _0516_ _3084_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3905_ _0564_ _0579_ _0600_ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__and4_1
X_6168__38 clknet_1_1__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__inv_2
X_4885_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] vssd1 vssd1 vccd1
+ vccd1 _1597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3836_ _2908_ _3093_ _0550_ _0552_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3767_ _2938_ _2926_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__nand2_1
X_5506_ _3002_ _0872_ _0420_ _0873_ _2211_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__a221oi_1
X_6486_ net60 _0319_ net46 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_3698_ _0417_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0418_
+ sky130_fd_sc_hd__nand2_1
X_5437_ _0941_ _0464_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5368_ _0835_ _0988_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4319_ _0816_ _2990_ _0817_ _2820_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__a221oi_1
X_5299_ _2005_ _2006_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__nor2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4670_ _0818_ _2824_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3621_ egd_top.BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__clkbuf_8
X_6340_ net82 _0173_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[90\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3552_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3483_ _2893_ _2985_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5222_ _1929_ _1930_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__nor2_1
X_5153_ _0378_ _0857_ _0341_ _0858_ _1861_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__a221oi_1
X_4104_ _0820_ _2810_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__nand2_1
X_5084_ _0992_ _2990_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4035_ _0397_ _0435_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _2560_ _2511_ _2557_ _2562_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__o211a_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4937_ _1647_ _0889_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 _2864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _0610_ _0922_ _0871_ _0921_ _1579_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_20 _1654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3819_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_42 egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4799_ _0650_ _0843_ _1510_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__o21ai_1
X_6469_ net211 _0302_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5840_ net16 _0920_ _2420_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__mux2_1
X_5771_ _2385_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4722_ _0881_ _3084_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4653_ _1365_ _1366_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__nand2_1
X_3604_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__buf_4
X_4584_ _2904_ _0872_ _0830_ _0873_ _1297_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__a221oi_1
X_3535_ _3083_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__buf_2
X_3466_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5205_ _0439_ _3048_ _0441_ _3002_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__a22o_1
X_3397_ _2883_ _2855_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__nor2_4
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5136_ _2914_ _0826_ _0506_ _0827_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__o22ai_1
X_5067_ _0602_ _3080_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__or2_1
X_4018_ _0357_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _0736_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5969_ _2495_ _2466_ _2545_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__nand3_1
Xclkbuf_0__2718_ _2718_ vssd1 vssd1 vccd1 vccd1 clknet_0__2718_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3320_ _2843_ egd_top.BitStream_buffer.pc\[2\] _2868_ vssd1 vssd1 vccd1 vccd1 _2869_
+ sky130_fd_sc_hd__and3_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__buf_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _2742_ _2748_ _2749_ _2751_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__o211ai_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823_ _2417_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ _2773_ _2774_ egd_top.BitStream_buffer.buffer_index\[4\] _2793_ vssd1 vssd1
+ vccd1 vccd1 _2376_ sky130_fd_sc_hd__or4b_4
XFILLER_0_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5685_ net4 _3112_ _2335_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4705_ _1417_ _0889_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4636_ _0990_ _0443_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4567_ _2867_ _3090_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nand2_1
X_4498_ _1211_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__nor2_1
X_3518_ _3066_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__inv_2
X_3449_ _2997_ _2812_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__nand2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _0538_ _0790_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__o21ai_1
X_6099_ _2667_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5470_ _2174_ _2175_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4421_ _0777_ _0781_ _2990_ _0782_ _1135_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4352_ _3008_ _0882_ _1064_ _1065_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__o2111a_1
X_4283_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__buf_4
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _2851_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__clkbuf_4
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _2505_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1
+ vccd1 _2597_ sky130_fd_sc_hd__nand2_1
X_3234_ net7 _2791_ _2798_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__mux2_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _2732_ _2733_ _0328_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout37 net38 vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3998_ _3123_ _2935_ _3126_ _0395_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__a22o_1
X_5806_ net36 egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__nand2_1
Xfanout48 net49 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
X_5737_ net10 _0463_ _2352_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5668_ _2329_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
X_4619_ _0937_ _0366_ _2957_ _0938_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__a221oi_1
X_5599_ net11 _0551_ _2281_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6189__58 clknet_1_0__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__inv_2
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _0992_ _3053_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__nand2_1
X_3921_ _2903_ _0638_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3852_ _3144_ _0335_ _3147_ _0338_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3783_ _2973_ _0333_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nand2_1
X_5522_ _3015_ _0987_ _2993_ _0989_ _2227_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5453_ _2153_ _2155_ _2157_ _2159_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4404_ _2881_ _0987_ _1116_ _0989_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__a221oi_2
X_5384_ _0865_ _2926_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4335_ _2959_ _2840_ _2847_ _0657_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__a221oi_2
X_4266_ _2922_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4197_ _3127_ _3096_ _3104_ _2859_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__a221oi_1
X_3217_ _2748_ _2746_ net30 vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__a21oi_1
X_6005_ _2577_ _2489_ _2580_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4120_ _0834_ _0836_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__nand2_1
X_4051_ _0434_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _0769_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 la_data_in_47_32[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4953_ _0407_ _3080_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3904_ _0605_ _0612_ _0617_ _0622_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4884_ _1594_ _1595_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3835_ _3104_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__nand2_1
X_3766_ _2934_ _0378_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6485_ net59 _0318_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_5505_ _2209_ _2210_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5436_ _0939_ _2939_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__nand2_1
X_3697_ _2933_ _2872_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5367_ _0833_ _2828_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__nand2_1
X_4318_ _1032_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5298_ _0567_ _0445_ _0686_ _0448_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__o22ai_1
X_4249_ _0435_ _0961_ _0962_ _0366_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3620_ _2899_ _2910_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3551_ _3099_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3482_ _3030_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__clkinv_4
X_6270_ clknet_1_0__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__buf_1
X_5221_ _0933_ _0610_ _0934_ _0443_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__a22o_1
X_5152_ _0337_ _2912_ _1403_ _2917_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__o22ai_1
X_4103_ _3004_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__clkbuf_4
X_5083_ _0990_ _3002_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4034_ _0394_ _0378_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5985_ _2479_ _2561_ _2512_ _2480_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__o211a_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_10 _0757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _0447_ _0923_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__o21ai_1
XANTENNA_32 _2927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _1724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_43 egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _2990_ _3055_ _3056_ _2808_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__a221oi_1
X_4798_ _0844_ _3002_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ _0463_ _2840_ _2847_ _0464_ _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__a221oi_2
X_6468_ net210 _0301_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_6399_ net141 _0232_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[57\]
+ sky130_fd_sc_hd__dfrtp_4
X_5419_ _3099_ _3017_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5770_ net15 _3030_ _2377_ vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4721_ _0516_ _3080_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4652_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] vssd1 vssd1 vccd1
+ vccd1 _1366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3603_ _2927_ _2985_ vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4583_ _1295_ _1296_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__nand2_1
X_6322_ clknet_1_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__buf_1
X_3534_ _2864_ _2871_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__nand2_1
X_3465_ _2899_ _2915_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__and2_1
X_5204_ _0464_ _0996_ _0657_ _0997_ _1912_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__a221oi_1
X_3396_ _2845_ _2872_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__nand2_1
X_5135_ _0816_ _2800_ _0817_ _0777_ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5066_ _2974_ _3096_ _3104_ _0657_ _1775_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _0722_ _0726_ _0729_ _0734_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5968_ _2543_ _2544_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__nand2_1
X_6224__90 clknet_1_1__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
XFILLER_0_47_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4919_ _3040_ _0848_ _2863_ _0849_ _1629_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2717_ _2717_ vssd1 vssd1 vccd1 vccd1 clknet_0__2717_ sky130_fd_sc_hd__clkbuf_16
X_5899_ _2474_ _2475_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _2809_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__clkbuf_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__inv_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5822_ net37 egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__nand2_1
X_5753_ _2375_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4704_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__inv_2
X_5684_ _2338_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4635_ _0981_ _0406_ _0982_ _3040_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4566_ _0841_ _0840_ _2881_ _0842_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__a221oi_1
X_3517_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__buf_4
X_4497_ _0933_ _0871_ _0934_ _0420_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__a22o_1
X_3448_ _2893_ _2996_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__and2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _2927_ _2769_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _0791_ _0330_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__nand2_1
X_6098_ _2665_ _2666_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__nand2_1
X_5049_ _0895_ _1011_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6203__71 clknet_1_1__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
XFILLER_0_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4420_ egd_top.BitStream_buffer.BS_buffer\[0\] _0783_ _0784_ _0625_ vssd1 vssd1 vccd1
+ vccd1 _1135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4351_ _1066_ _0889_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__or2_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _0432_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__clkbuf_4
X_3302_ _2850_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__inv_2
X_3233_ _2797_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__buf_4
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _2516_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1
+ vccd1 _2596_ sky130_fd_sc_hd__nand2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _2736_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout38 net46 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3997_ _0561_ _3110_ _0712_ _0713_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__o2111a_1
X_5805_ _2406_ _2408_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[5\] sky130_fd_sc_hd__nor2_2
Xfanout49 net50 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_4
X_5736_ _2365_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5667_ net11 _0336_ _2317_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__mux2_1
X_4618_ _1330_ _1331_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5598_ _2292_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
X_4549_ _1252_ _1255_ _1258_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__and4_1
X_6273__135 clknet_1_1__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3920_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__buf_4
X_3851_ _0568_ _0569_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3782_ _2971_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _0501_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5521_ _2225_ _2226_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5452_ _0974_ _3112_ _0975_ _3119_ _2158_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__a221oi_1
X_4403_ _1117_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nand2_1
X_5383_ _2081_ _2084_ _2087_ _2089_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__and4_1
X_4334_ _0619_ _2854_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4265_ _0413_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__clkbuf_4
X_6004_ _2578_ _2579_ _2500_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__o21ai_1
X_4196_ _0641_ _3093_ _0912_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__o21ai_1
X_3216_ _2784_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6194__62 clknet_1_0__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__inv_2
X_5719_ net4 _0435_ _2353_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__2731_ clknet_0__2731_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2731_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4050_ _0432_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0768_
+ sky130_fd_sc_hd__nand2_1
Xinput6 la_data_in_47_32[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_4
XFILLER_0_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _0343_ _3096_ _3104_ _0495_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3903_ _0618_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__nor2_1
X_4883_ _1116_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3834_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__clkbuf_8
X_6304__164 clknet_1_1__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__inv_2
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3765_ _0468_ _0473_ _0479_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and4_1
X_6484_ net58 _0317_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_6325__15 clknet_1_1__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__inv_2
X_5504_ _0877_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _2210_
+ sky130_fd_sc_hd__nand2_1
X_3696_ _0410_ _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__nor2_1
X_5435_ _0638_ _0921_ _3002_ _0922_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5366_ _0824_ _0395_ _0825_ _2935_ _2072_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4317_ _0820_ _2812_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5297_ _0438_ _3002_ _0440_ _3030_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__a22o_1
X_4248_ _3133_ _0963_ _0575_ _0964_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__o22ai_1
X_4179_ _0895_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _0896_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6279__141 clknet_1_0__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _2856_ _2871_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6173__43 clknet_1_0__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__inv_2
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3481_ egd_top.BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__clkbuf_8
X_5220_ egd_top.BitStream_buffer.BS_buffer\[77\] _0930_ _0931_ egd_top.BitStream_buffer.BS_buffer\[80\]
+ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__a22o_1
X_5151_ _0920_ _2840_ _2847_ _0587_ _1859_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__a221oi_1
X_4102_ _0818_ _2816_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__nand2_1
X_5082_ _0981_ _0402_ _0982_ _2863_ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__a221oi_1
X_4033_ _0391_ _3139_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5984_ _2466_ _2488_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4935_ _0885_ _3101_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 _0757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _0925_ _0583_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__nand2_1
XANTENNA_22 _1767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4797_ _1498_ _1502_ _1504_ _1508_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__and4_1
XANTENNA_44 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 _2927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _0534_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__nand2_1
X_3748_ _0465_ _2854_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3679_ _0397_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6467_ net209 _0300_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_6398_ net140 _0231_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_5418_ _3139_ _0907_ _3105_ _0908_ _2124_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__a221oi_1
X_5349_ _2808_ _0787_ _3124_ _0788_ _2055_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4720_ _0378_ _3096_ _3104_ _0464_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4651_ _1363_ _1364_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3602_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4582_ _0877_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1296_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3533_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__inv_2
X_3464_ _3008_ _3009_ _3011_ _3012_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5203_ _1910_ _1911_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__nand2_1
X_5134_ _1841_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__nand2_1
X_3395_ _2943_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5065_ _0334_ _3093_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__o21ai_1
X_4016_ _0732_ _0733_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5967_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4918_ _0489_ _0850_ _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__o21ai_1
X_5898_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4849_ _0970_ _0976_ _0574_ _0977_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ net28 _2745_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5821_ _2762_ _2397_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[1\] sky130_fd_sc_hd__xor2_4
X_5752_ _2374_ _2794_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4703_ _0885_ _1116_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5683_ net5 _0346_ _2335_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4634_ _0506_ _0405_ _0756_ _0409_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__o22ai_1
X_4565_ _2944_ _0843_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__o21ai_1
X_3516_ _2927_ _2996_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__nand2_4
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4496_ egd_top.BitStream_buffer.BS_buffer\[71\] _0930_ _0931_ _2859_ vssd1 vssd1
+ vccd1 vccd1 _1211_ sky130_fd_sc_hd__a22o_1
X_3447_ _2961_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__buf_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ clknet_1_0__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__buf_1
X_3378_ _2883_ _2842_ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__nor2_8
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _2505_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1
+ vccd1 _2666_ sky130_fd_sc_hd__nand2_1
X_5117_ _2791_ _0782_ _1116_ _0781_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__a221oi_2
X_5048_ _0443_ _0872_ _0587_ _0873_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6250__114 clknet_1_1__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__inv_2
X_3301_ egd_top.BitStream_buffer.pc\[5\] _2768_ _2834_ vssd1 vssd1 vccd1 vccd1 _2850_
+ sky130_fd_sc_hd__or3_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ _0428_ _2959_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__nand2_1
X_3232_ _2796_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__buf_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _2519_ _2526_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__nor2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _2734_ _2735_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5804_ _2405_ _2394_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3996_ _3118_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _0714_
+ sky130_fd_sc_hd__nand2_1
Xfanout39 net41 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_4
XFILLER_0_91_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5735_ net11 _2830_ _2353_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5666_ _2328_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4617_ _0941_ _3105_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5597_ net12 _3101_ _2281_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__mux2_1
X_4548_ _0330_ _0800_ _0801_ _2818_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__a221oi_1
X_4479_ _2952_ _3131_ _0347_ _3135_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__o22ai_1
X_6218_ clknet_1_1__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__buf_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _2714_ _2715_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__nand2_1
XFILLER_0_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _2800_ _3157_ _0329_ _2791_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3781_ _2969_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0500_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5520_ _0992_ _3070_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5451_ _0543_ _0976_ _3129_ _0977_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__o22ai_1
X_4402_ _0992_ _3034_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__nand2_1
X_5382_ _0343_ _0857_ _2974_ _0858_ _2088_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4333_ _2858_ _0464_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__nand2_1
X_4264_ _0411_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3215_ _2747_ net30 _2783_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__mux2_1
X_6003_ _2454_ _2531_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__nor2_1
X_4195_ _3100_ _2943_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5718_ _2356_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_1
X_3979_ _3058_ _3055_ _3056_ _2810_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ net5 _3124_ _2317_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__2730_ clknet_0__2730_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2730_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6256__120 clknet_1_1__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
Xinput7 la_data_in_47_32[15] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
X_6318__9 clknet_1_0__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__inv_2
X_4951_ _1519_ _3093_ _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3902_ _0619_ _0446_ _0620_ _0449_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _1541_ _0903_ _1593_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3833_ _3100_ _0551_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3764_ _0481_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6483_ net57 _0316_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_3695_ _0411_ _0412_ _0413_ _0414_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__a22o_1
X_5503_ _0874_ _0443_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__nand2_1
X_5434_ _0444_ _0923_ _2140_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5365_ _0506_ _0826_ _2908_ _0827_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4316_ _0818_ _2818_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__nand2_1
X_5296_ egd_top.BitStream_buffer.BS_buffer\[79\] _0996_ egd_top.BitStream_buffer.BS_buffer\[82\]
+ _0997_ _2003_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__a221oi_2
X_4247_ _3148_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__clkbuf_4
X_4178_ _2962_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__clkbuf_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3480_ _2995_ _3006_ _3019_ _3028_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5150_ _0789_ _2854_ _1858_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__o21ai_1
X_4101_ _2999_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__clkbuf_4
X_5081_ _0641_ _0405_ _0506_ _0409_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4032_ _0388_ _0392_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5983_ _2558_ _2559_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4934_ _0883_ _0551_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _0772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _1565_ _1569_ _1573_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__and4_1
XANTENNA_23 _2064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4796_ _0742_ _0831_ _0832_ _2824_ _1507_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__a221oi_2
XANTENNA_45 _0583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_34 _2946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ _3060_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _0535_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3747_ _2858_ _2830_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3678_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__buf_4
X_6466_ net208 _0299_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6397_ net139 _0230_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5417_ _1417_ _3109_ _2123_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__o21ai_1
X_5348_ _0795_ _0790_ _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__o21ai_1
X_5279_ _1985_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4650_ _0469_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3601_ _3139_ _3141_ _2771_ _3142_ _3149_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__a221oi_1
Xinput10 la_data_in_47_32[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4581_ _0874_ _0583_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__nand2_1
X_3532_ _3078_ _3080_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__or2_1
X_3463_ _2895_ _2915_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5202_ _0999_ _0871_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__nand2_1
X_5133_ _0820_ _2826_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__nand2_1
X_3394_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ _3100_ _0406_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4015_ _0352_ egd_top.BitStream_buffer.BS_buffer\[0\] _0353_ egd_top.BitStream_buffer.BS_buffer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _2542_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5897_ _2473_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4917_ _2867_ _3124_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4848_ _0967_ _0469_ _0968_ _0988_ _1559_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4779_ _0802_ _2804_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6449_ net191 _0282_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5820_ _2416_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5751_ egd_top.BitStream_buffer.buffer_index\[4\] net224 vssd1 vssd1 vccd1 vccd1
+ _2374_ sky130_fd_sc_hd__or2_1
X_4702_ _0883_ _0841_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5682_ _2337_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4633_ _1340_ _1342_ _1344_ _1346_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4564_ _0844_ _3034_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__nand2_1
X_3515_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4495_ _0587_ _0921_ _2904_ _0922_ _1209_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__a221oi_1
X_3446_ _2981_ _2982_ _2988_ _2991_ _2994_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _2516_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] vssd1 vssd1 vccd1
+ vccd1 _2665_ sky130_fd_sc_hd__nand2_1
X_5116_ egd_top.BitStream_buffer.BS_buffer\[6\] _0783_ _0784_ _0988_ vssd1 vssd1 vccd1
+ vccd1 _1825_ sky130_fd_sc_hd__a22o_1
X_5047_ _1755_ _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5949_ _2524_ _2525_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3300_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ _0430_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3231_ _2773_ _2795_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__or2_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ net33 net32 vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5803_ _2407_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3995_ _3114_ _0389_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__nand2_1
X_5734_ _2364_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
X_5665_ net12 _3143_ _2317_ vssd1 vssd1 vccd1 vccd1 _2328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4616_ _0939_ _0333_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5596_ _2291_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
X_4547_ _1259_ _1260_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4478_ _1147_ _1161_ _1174_ _1192_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__and4_1
X_3429_ _2970_ _2972_ _2975_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__and4_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _2691_ _2702_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__nand2_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _2646_ _2648_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3780_ _2956_ _0371_ _2958_ _0495_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5450_ _0967_ _0551_ _0968_ _2881_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4401_ _0990_ _0638_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5381_ _3133_ _2911_ _0334_ _2916_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4332_ _2887_ _0848_ _0406_ _0849_ _1047_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__a221oi_1
X_4263_ _0960_ _0966_ _0973_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3214_ _2781_ _2782_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__nand2_1
X_6002_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _2532_ vssd1 vssd1
+ vccd1 vccd1 _2578_ sky130_fd_sc_hd__nor2_1
X_4194_ egd_top.BitStream_buffer.BS_buffer\[54\] _0907_ _2951_ _0908_ _0910_ vssd1
+ vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _0694_ _0695_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__nand2_1
X_5717_ net5 _0366_ _2353_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5648_ _2319_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5579_ net6 _0625_ _2281_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 la_data_in_47_32[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4950_ _3100_ _3010_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__nand2_1
X_3901_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__inv_2
X_4881_ _1554_ _1563_ _1577_ _1592_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and4_1
X_3832_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5502_ _3142_ _0863_ _0864_ _2951_ _2207_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__a221oi_2
X_3763_ _2919_ _2922_ _2921_ _2913_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6482_ net56 _0315_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[117\]
+ sky130_fd_sc_hd__dfrtp_1
X_3694_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5433_ _0925_ _0477_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__nand2_1
X_5364_ _0816_ _2804_ _0817_ _0886_ _2070_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__a221oi_1
X_4315_ _3030_ _0809_ _3070_ _0810_ _1030_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5295_ _2001_ _2002_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__nand2_1
X_4246_ _3145_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__clkbuf_4
X_4177_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__buf_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6286__147 clknet_1_0__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__inv_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6330__20 clknet_1_0__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__inv_2
X_4100_ _2997_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__clkbuf_4
X_5080_ _1783_ _1785_ _1787_ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__and4_1
X_4031_ _0745_ _0746_ _0747_ _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5982_ egd_top.exp_golomb_decoding.te_range\[2\] vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4933_ _0610_ _0872_ _0875_ _0873_ _1643_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__a221oi_1
Xclkbuf_0__2731_ _2731_ vssd1 vssd1 vccd1 vccd1 clknet_0__2731_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4864_ _1574_ _1575_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__nor2_1
XANTENNA_13 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _1505_ _1506_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__nand2_1
XANTENNA_24 _2160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 _2816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _2979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3815_ _3057_ _3066_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__nand2_1
X_3746_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6465_ net207 _0298_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3677_ _2927_ _2837_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5416_ _3117_ _0398_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__nand2_1
X_6396_ net138 _0229_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_5347_ _0791_ _2800_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _0897_ _0830_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__nand2_1
X_4229_ _0377_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3600_ _3144_ _3145_ _3147_ _3148_ vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__o22ai_1
Xinput11 la_data_in_47_32[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_4
X_4580_ egd_top.BitStream_buffer.BS_buffer\[55\] _0863_ _0864_ egd_top.BitStream_buffer.BS_buffer\[53\]
+ _1293_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3531_ _3079_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__buf_2
XFILLER_0_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3462_ _3010_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5201_ _0428_ _0875_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__nand2_1
X_3393_ _2926_ _2929_ _2930_ _2931_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__a221oi_2
X_5132_ _0818_ _0625_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _2951_ _0907_ _2957_ _0908_ _1772_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4014_ _0730_ _0348_ _0731_ _0350_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5965_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5896_ _2463_ _2789_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4916_ _2881_ _0840_ _0414_ _0842_ _1626_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__a221oi_1
X_4847_ _0717_ _0969_ _0543_ _0971_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4778_ _1488_ _3065_ _0795_ _0796_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3729_ _0448_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__buf_4
XFILLER_0_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6448_ net190 _0281_ net42 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_6379_ net121 _0212_ net51 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[77\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6215__82 clknet_1_0__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6230__96 clknet_1_1__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5750_ _2373_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
X_5681_ net6 _2926_ _2335_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4701_ _0477_ _0872_ _0926_ _0873_ _1413_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__a221oi_1
X_4632_ _0974_ _3146_ _0975_ _3132_ _1345_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4563_ _1266_ _1270_ _1272_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3514_ _3053_ _3055_ _3056_ _2806_ _3062_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__a221oi_1
X_4494_ _1207_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__nand2_1
X_3445_ _2992_ _2993_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__nand2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _2862_ _2890_ _2906_ _2924_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__and4_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _2595_ _2663_ _2635_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__nand3_1
X_5115_ _1823_ _1824_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__nand2_1
X_5046_ _0877_ _0346_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5948_ _2505_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1
+ vccd1 _2525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5879_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] _2455_ vssd1 vssd1
+ vccd1 vccd1 _2456_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _2774_ _2794_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__or2_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _2732_ _2733_ _2734_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5802_ net35 egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__nand2_1
X_3994_ _3111_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _0712_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5733_ net12 _2859_ _2353_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5664_ _2327_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
X_4615_ _1327_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5595_ net13 _0841_ _2281_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__mux2_1
X_4546_ _0804_ _2826_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4477_ _1178_ _1182_ _1187_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__and4_1
X_3428_ _2976_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _2977_
+ sky130_fd_sc_hd__nand2_1
X_3359_ _2907_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__inv_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _2711_ _2554_ _2713_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__nand3_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _2616_ _2647_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__nand2_2
X_5029_ _0844_ _3037_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4400_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5380_ _0587_ _2839_ _2846_ _0583_ _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__a221oi_1
X_4331_ _3082_ _0850_ _1046_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__o21ai_1
X_4262_ _0974_ _0333_ _0975_ _3143_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3213_ _2732_ _2739_ net34 net32 vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__and4_1
X_6001_ _2576_ _2469_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4193_ _0717_ _3110_ _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3977_ _3060_ _2818_ vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5716_ _2355_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5647_ net6 _3127_ _2317_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__mux2_1
X_5578_ _2282_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__clkbuf_1
X_4529_ _1242_ _1243_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__nor2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6185__54 clknet_1_0__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__inv_2
XFILLER_0_36_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 la_data_in_47_32[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6263__126 clknet_1_1__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4880_ _1580_ _1584_ _1588_ _1591_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__and4_1
X_3900_ _2987_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__clkinv_4
X_3831_ _3096_ _3090_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3762_ _0480_ _2912_ _2981_ _2917_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o22ai_1
X_5501_ _2205_ _2206_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6481_ net55 _0314_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_3693_ _2767_ _2872_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__and2_1
X_5432_ _2987_ _0933_ _3034_ _0934_ _2138_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5363_ _2068_ _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__nand2_1
X_4314_ _0480_ _0811_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5294_ _0999_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _2002_
+ sky130_fd_sc_hd__nand2_1
X_4245_ _2771_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4176_ _2958_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _0384_ _2951_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5981_ net21 _2557_ net20 vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__and3b_1
X_4932_ _1641_ _1642_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2730_ _2730_ vssd1 vssd1 vccd1 vccd1 clknet_0__2730_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4863_ _0789_ _0446_ _1005_ _0449_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__o22ai_1
XANTENNA_14 _0841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4794_ _0835_ _0777_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__nand2_1
XANTENNA_25 _2162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _0531_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__nor2_1
XANTENNA_36 _3031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__clkbuf_8
X_6164__35 clknet_1_1__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__inv_2
XFILLER_0_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6464_ net206 _0297_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6310__1 clknet_1_1__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__inv_2
X_3676_ _0394_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__nand2_1
X_5415_ _2110_ _2114_ _2118_ _2121_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6395_ net137 _0228_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_5346_ _2802_ _0782_ _3101_ _0781_ _2052_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5277_ _0895_ _2874_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__nand2_1
X_4228_ _0380_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__clkbuf_4
X_4159_ _0874_ _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__nand2_1
X_6246__110 clknet_1_1__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 la_data_in_47_32[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3530_ _2833_ _2871_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3461_ egd_top.BitStream_buffer.BS_buffer\[19\] vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__buf_4
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5200_ _3010_ _0987_ _0414_ _0989_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__a221oi_1
X_3392_ _2936_ _2940_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__nand2_1
X_5131_ _2808_ _0810_ _3070_ _0809_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5062_ _1066_ _3110_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__o21ai_1
X_4013_ _2939_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6269__132 clknet_1_0__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5964_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5895_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] _2470_ _2471_ vssd1
+ vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__o21ai_1
X_4915_ _0881_ _0843_ _1625_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__o21ai_1
X_4846_ _0553_ _0961_ _0962_ _3105_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _0797_ _2810_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__nand2_1
X_3728_ _2845_ _2852_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__nand2_1
X_3659_ _0377_ _0378_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__nand2_1
X_6447_ net189 _0280_ net38 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_6378_ net120 _0211_ net51 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[78\]
+ sky130_fd_sc_hd__dfrtp_4
X_5329_ _2025_ _2028_ _2032_ _2036_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5680_ _2336_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
X_4700_ _1411_ _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nand2_1
X_4631_ _0575_ _0976_ _0970_ _0977_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4562_ _0875_ _0831_ _0832_ _2820_ _1275_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__a221oi_1
X_3513_ _3059_ _3061_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__nand2_1
X_4493_ _0925_ _0875_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3444_ egd_top.BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__buf_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3375_ _2918_ _2923_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__nor2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _2573_ _2598_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__nor2_1
X_5114_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1
+ vccd1 _1824_ sky130_fd_sc_hd__nand2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _0874_ _2904_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5947_ _2516_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1
+ vccd1 _2524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5878_ _2453_ _2454_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__nand2_1
X_4829_ _1495_ _1509_ _1522_ _1540_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ net222 vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__inv_2
Xhold1 net225 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ egd_top.BitStream_buffer.pc_reg\[6\] _2406_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[6\]
+ sky130_fd_sc_hd__xor2_4
X_3993_ _0480_ _3093_ _0707_ _0708_ _0710_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__o2111a_1
X_5732_ _2363_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ net13 _0333_ _2317_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4614_ _0933_ _0420_ _0934_ _0607_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5594_ _2290_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
X_4545_ _0802_ _2800_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4476_ _0892_ _0709_ _0893_ _0830_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__a221oi_1
X_3427_ _2964_ _2852_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__and2_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _2712_ _2514_ _2705_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__nand3_1
X_3358_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__buf_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _2555_ _2589_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__nor2_1
X_3289_ _2833_ _2837_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__and2_1
X_5028_ _1727_ _1731_ _1733_ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4330_ _2867_ _2980_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__nand2_1
X_4261_ _3147_ _0976_ _0349_ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__o22ai_1
X_3212_ _2742_ _2748_ _2752_ _2778_ _2780_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__o2111ai_1
X_6000_ _2447_ _2467_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4192_ _3118_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _0909_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2719_ clknet_0__2719_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2719_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6240__105 clknet_1_1__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XFILLER_0_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3976_ _3057_ _3153_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5715_ net6 _0398_ _2353_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5646_ _2318_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5577_ net7 _0458_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4528_ _3031_ _0446_ _0444_ _0449_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__o22ai_1
X_4459_ _1164_ _1167_ _1170_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__and4_1
X_6129_ _2674_ _2512_ _2645_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__nand3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3830_ _0543_ _3077_ _0545_ _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__o2111a_1
X_3761_ _3127_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__inv_2
X_5500_ _0867_ _0392_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6480_ net54 _0313_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3692_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5431_ egd_top.BitStream_buffer.BS_buffer\[79\] _0930_ _0931_ _0894_ vssd1 vssd1
+ vccd1 vccd1 _2138_ sky130_fd_sc_hd__a22o_1
X_5362_ _0820_ _0458_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__nand2_1
X_4313_ _0812_ _3015_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nand2_1
X_5293_ _0427_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _2001_
+ sky130_fd_sc_hd__nand2_1
X_4244_ _3141_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__clkbuf_4
X_4175_ _2956_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3959_ _3011_ _3009_ _0602_ _3012_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__o22ai_1
X_5629_ net13 _2863_ _2299_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5980_ _2556_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4931_ _0877_ _2926_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4862_ _0439_ _0443_ _0441_ _2987_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3813_ _3047_ _3002_ egd_top.BitStream_buffer.BS_buffer\[126\] _3050_ vssd1 vssd1
+ vccd1 vccd1 _0532_ sky130_fd_sc_hd__a22o_1
X_4793_ _0833_ _2818_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__nand2_1
XANTENNA_37 _3078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 _2902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_26 _2276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 _0886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3744_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3675_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6463_ net205 _0296_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5414_ _2119_ _2120_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6394_ net136 _0227_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_5345_ _1116_ _0783_ _0784_ _0841_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5276_ _3034_ _0872_ _0583_ _0873_ _1983_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__a221oi_1
X_4227_ _0937_ _3142_ _0398_ _0938_ _0943_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__a221oi_2
X_4158_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4089_ _0803_ _0805_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6292__153 clknet_1_1__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__inv_2
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput13 la_data_in_47_32[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_4
X_3460_ _2927_ _2915_ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__nand2_1
X_3391_ _2938_ _2939_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__nand2_1
X_5130_ _1519_ _0811_ _1838_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5061_ _3118_ _0392_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__nand2_1
X_4012_ _3119_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5963_ _2537_ _2539_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4914_ _0844_ _3030_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5894_ _2459_ _2451_ _2449_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__and3_1
X_4845_ _0347_ _0963_ _0730_ _0964_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__o22ai_1
X_4776_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__inv_2
X_3727_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3658_ egd_top.BitStream_buffer.BS_buffer\[37\] vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6446_ net188 _0279_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3589_ _3089_ _3107_ _3121_ _3137_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__and4_1
X_6377_ net119 _0210_ net51 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[79\]
+ sky130_fd_sc_hd__dfrtp_4
X_5328_ _0926_ _0945_ _0946_ _2926_ _2035_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__a221oi_1
X_5259_ _0414_ _0840_ _2993_ _0842_ _1966_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__a221oi_1
X_6300__160 clknet_1_0__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__inv_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6206__73 clknet_1_0__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4630_ _0967_ _0886_ _0968_ _2874_ _1343_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__a221oi_1
X_6221__87 clknet_1_0__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
XFILLER_0_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6299__159 clknet_1_0__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__inv_2
XFILLER_0_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4561_ _1273_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3512_ _3060_ _2814_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__nand2_1
X_4492_ _0923_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _1207_
+ sky130_fd_sc_hd__or2b_1
X_6231_ clknet_1_1__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__buf_1
X_3443_ _2946_ _2915_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__and2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _1821_ _1822_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__nand2_1
X_3374_ _2919_ _2920_ _2921_ _2922_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__a22o_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _2660_ _2661_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__nand2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _0385_ _0863_ _0864_ egd_top.BitStream_buffer.BS_buffer\[57\] _1753_ vssd1
+ vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5946_ _2519_ _2522_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5877_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] vssd1 vssd1 vccd1 vccd1
+ _2454_ sky130_fd_sc_hd__inv_4
XFILLER_0_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4828_ _1526_ _1530_ _1535_ _1539_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4759_ _1470_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6429_ net171 _0262_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 net34 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3992_ _3104_ _0709_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nand2_1
X_5800_ _2394_ _2405_ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5731_ net13 _0709_ _2353_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5662_ _2326_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
X_4613_ egd_top.BitStream_buffer.BS_buffer\[72\] _0930_ _0931_ egd_top.BitStream_buffer.BS_buffer\[75\]
+ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__a22o_1
X_5593_ net14 _1116_ _2281_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__mux2_1
X_4544_ _1256_ _3065_ _0538_ _0796_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__o221a_1
X_4475_ _1188_ _1189_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__nand2_1
X_3426_ _2973_ _2974_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__nand2_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _2697_ _2691_ _2651_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3357_ _2891_ _2894_ _2897_ _2901_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__o2111a_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _2645_ _2512_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__nand2_1
X_5027_ _0871_ _0831_ _0832_ _2828_ _1736_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__a221oi_1
X_3288_ _2836_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5929_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1 vccd1
+ _2506_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6200__68 clknet_1_1__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__inv_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4260_ _0338_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4191_ _3114_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__buf_4
X_3211_ egd_top.BitStream_buffer.pc\[6\] _2751_ _2771_ _2779_ vssd1 vssd1 vccd1 vccd1
+ _2780_ sky130_fd_sc_hd__or4b_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2718_ clknet_0__2718_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2718_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3975_ _0691_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5714_ _2354_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
X_5645_ net7 _2907_ _2317_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5576_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4527_ _0439_ egd_top.BitStream_buffer.BS_buffer\[95\] _0441_ _0638_ vssd1 vssd1
+ vccd1 vccd1 _1242_ sky130_fd_sc_hd__a22o_1
X_4458_ _3090_ _0857_ _2907_ _0858_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__a221oi_1
X_3409_ _2767_ _2837_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__and2_1
X_4389_ _1005_ _0956_ _3064_ _0958_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o22ai_2
X_6128_ _2649_ _2691_ _2677_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__nand3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _2630_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3760_ _0474_ _2894_ _0475_ _0476_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_27_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3691_ _2902_ _2872_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__and2_1
X_5430_ _2122_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _0818_ _1011_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4312_ _1016_ _1020_ _1023_ _1027_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5292_ _0406_ _0987_ _2887_ _0989_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__a221oi_1
X_4243_ _2804_ _0954_ _2802_ _0955_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__a221oi_2
X_4174_ _0881_ _0882_ _0884_ _0887_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3958_ _0672_ _0673_ _0674_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__and4_1
XFILLER_0_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3889_ _0419_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5628_ _2308_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5559_ _2253_ _2256_ _2260_ _2264_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4930_ _0874_ _0607_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4861_ _2830_ _0996_ _0464_ _0997_ _1572_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_47_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3812_ egd_top.BitStream_buffer.BS_buffer\[124\] _3043_ _3044_ egd_top.BitStream_buffer.BS_buffer\[125\]
+ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__a22o_1
X_4792_ _0824_ _3097_ _0825_ _3090_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__a221oi_1
XANTENNA_38 _3078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _2771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 _0988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_49 _2927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3743_ _0460_ _0462_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__nand2_1
X_3674_ _2895_ _2909_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__and2_1
X_6462_ net204 _0295_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6393_ net135 _0226_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_5413_ _0723_ _0445_ _0789_ _0448_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5344_ _2050_ _2051_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__nand2_1
X_6321__12 clknet_1_0__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__inv_2
XFILLER_0_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5275_ _1981_ _1982_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__nand2_1
X_4226_ _0940_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4157_ _2969_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__clkbuf_4
X_4088_ _0804_ _2820_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__nand2_1
X_6227__93 clknet_1_1__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
XFILLER_0_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6155__26 clknet_1_0__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__inv_2
XFILLER_0_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 la_data_in_47_32[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
XFILLER_0_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3390_ egd_top.BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5060_ _0336_ _3126_ _3146_ _3123_ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__a221oi_1
X_4011_ _0727_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _2468_ _2538_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4913_ _1613_ _1617_ _1619_ _1623_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5893_ _2469_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4844_ _2814_ _0954_ _2812_ _0955_ _1555_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4775_ _2791_ _0787_ _2980_ _0788_ _1486_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3726_ _0445_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__clkbuf_4
X_6276__138 clknet_1_0__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
X_3657_ _2870_ _2910_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__and2_1
X_6445_ net187 _0278_ net44 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3588_ _3128_ _3136_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__nor2_1
X_6376_ net118 _0209_ net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5327_ _2033_ _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__nand2_1
X_5258_ _3011_ _0843_ _1965_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__o21ai_1
X_5189_ _2830_ _0961_ _0962_ _2859_ _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__a221oi_1
X_4209_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ _0835_ _0458_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4491_ _1195_ _1198_ _1201_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__and4_1
X_3511_ _2964_ _2961_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__and2_1
X_3442_ _2989_ _2990_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__nand2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__buf_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5112_ _3101_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _2656_ _2513_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__nand2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _1751_ _1752_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5945_ _2520_ _2521_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__nand2_1
X_5876_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1 vccd1 vccd1
+ _2453_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4827_ _0892_ _0463_ _0893_ _0875_ _1538_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758_ _0999_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _1471_
+ sky130_fd_sc_hd__nand2_1
X_3709_ _0428_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _0429_
+ sky130_fd_sc_hd__nand2_1
X_4689_ _0894_ _2840_ _2847_ _0830_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__a221oi_1
X_6428_ net170 _0261_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6359_ net101 _0192_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6259__122 clknet_1_1__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 _2792_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3991_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5730_ _2362_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6307__167 clknet_1_1__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__inv_2
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5661_ net14 _2974_ _2317_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4612_ _0742_ _0921_ _0477_ _0922_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__a221oi_1
X_5592_ _2289_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
X_4543_ _0797_ _2806_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4474_ _0897_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _1189_
+ sky130_fd_sc_hd__nand2_1
X_3425_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__clkbuf_8
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _2710_ _2513_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__nand2_1
X_3356_ _2903_ _2904_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__nand2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _2639_ _2644_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__nand2_1
X_3287_ _2834_ _2835_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2836_
+ sky130_fd_sc_hd__and3_2
X_5026_ _1734_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__nand2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5928_ _2481_ _2499_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__nor2_4
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6197__65 clknet_1_0__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__inv_2
X_5859_ _2436_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3210_ _2774_ _2775_ egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1
+ vccd1 _2779_ sky130_fd_sc_hd__and3_1
X_4190_ _3111_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2717_ clknet_0__2717_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2717_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _3047_ _3030_ egd_top.BitStream_buffer.BS_buffer\[127\] _3050_ vssd1 vssd1
+ vccd1 vccd1 _0692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5713_ net7 _3139_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6328__18 clknet_1_1__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__inv_2
X_5644_ _2316_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5575_ _2793_ _2776_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__nand2_2
X_4526_ _0553_ _0996_ _2830_ _0997_ _1240_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__a221oi_1
X_4457_ _1171_ _2912_ _0480_ _2917_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3408_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__clkbuf_8
X_6127_ _2692_ _2513_ _2694_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4388_ _1092_ _1095_ _1099_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__and4_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _2886_ _2887_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__nand2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _2615_ _2560_ _2466_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__or3_1
X_5009_ _1717_ _3065_ _1140_ _0796_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6176__46 clknet_1_0__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__inv_2
X_3690_ _0403_ _0405_ _0407_ _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5360_ _2791_ _0809_ _2812_ _0810_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__a221oi_1
X_4311_ _3153_ _0800_ _0801_ _2814_ _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__a221oi_1
X_5291_ _1997_ _1998_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4242_ _0772_ _0956_ _0957_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__o22ai_1
X_4173_ _0888_ _0889_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__or2_1
X_3957_ _3004_ _2808_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3888_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__buf_8
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5627_ net14 _0402_ _2299_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5558_ _0875_ _0945_ _0946_ _3112_ _2263_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__a221oi_1
X_4509_ _2808_ _0954_ _2806_ _0955_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5489_ _3007_ _0840_ _0406_ _0842_ _2194_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4860_ _1570_ _1571_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__nand2_1
X_3811_ _0526_ _3032_ _0527_ _0528_ _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__o2111a_1
XANTENNA_39 _3082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4791_ _0601_ _0826_ _0983_ _0827_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__o22ai_1
XANTENNA_28 _2771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_17 _1192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3742_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] vssd1 vssd1
+ vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3673_ _0391_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__nand2_1
X_6461_ net203 _0294_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_6392_ net134 _0225_ net48 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_5412_ _0438_ _3030_ _0440_ _3037_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5343_ net221 egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1
+ vccd1 _2051_ sky130_fd_sc_hd__nand2_1
X_5274_ _0877_ _3119_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__nand2_1
X_4225_ _0941_ _2957_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__nand2_1
X_4156_ _2971_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4087_ _3060_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__clkbuf_4
X_4989_ _0941_ _2859_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6253__117 clknet_1_0__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 la_data_in_47_32[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
XFILLER_0_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4010_ _0340_ _2974_ _0342_ _0333_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a22o_1
X_5961_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4912_ _0583_ _0831_ _0832_ _2826_ _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_87_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5892_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] _2468_ vssd1 vssd1 vccd1
+ vccd1 _2469_ sky130_fd_sc_hd__nor2_1
X_4843_ _0686_ _0956_ _1021_ _0958_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _0723_ _0790_ _1485_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3725_ _2946_ _2984_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6444_ net186 _0277_ net46 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3656_ _0372_ _0375_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3587_ _3129_ _3131_ _3133_ _3135_ vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__o22ai_1
X_6375_ net117 _0208_ net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5326_ _0949_ _3105_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5257_ _0844_ _2990_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__nand2_1
X_4208_ _0359_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__clkbuf_4
X_5188_ _3075_ _0963_ _3108_ _0964_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__o22ai_1
X_4139_ _0464_ _2840_ _2847_ _0495_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3510_ _3057_ _3058_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4490_ _0717_ _3077_ _1202_ _1203_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__o2111a_1
X_6236__101 clknet_1_0__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
X_3441_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _2833_ _2915_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__and2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _1768_ _0903_ _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__nand3_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _2646_ _2648_ _2514_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__o21ai_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _0867_ _3115_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5944_ _2505_ _2437_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5875_ _2450_ _2451_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__nand2_1
X_4826_ _1536_ _1537_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4757_ _0428_ _1000_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3708_ _0427_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__buf_4
X_4688_ _1126_ _2854_ _1400_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__o21ai_1
X_6427_ net169 _0260_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_3639_ _2946_ _2852_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__and2_1
X_6358_ net100 _0191_ net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5309_ _3086_ _0366_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 _2793_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ _3100_ _2881_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5660_ _2325_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4611_ _1323_ _1324_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5591_ net15 _0988_ _2281_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__mux2_1
X_4542_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__inv_2
X_4473_ _0895_ _2826_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nand2_1
X_3424_ _2964_ _2909_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__buf_8
X_6143_ _2707_ _2709_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__nand2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6074_ _2641_ _2642_ _2496_ _2489_ _2643_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__o32a_1
X_3286_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__inv_2
X_5025_ _0835_ _0886_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__nand2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5927_ _2481_ _2499_ _2439_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ net1 _0477_ _2419_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5789_ egd_top.BitStream_buffer.pc_reg\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__or2_1
X_4809_ _3124_ _0857_ _0395_ _0858_ _1520_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5712_ _2352_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__buf_4
X_3973_ egd_top.BitStream_buffer.BS_buffer\[125\] _3043_ _3044_ egd_top.BitStream_buffer.BS_buffer\[126\]
+ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__a22o_1
X_6313__4 clknet_1_1__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__inv_2
XFILLER_0_17_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5643_ egd_top.BitStream_buffer.buffer_index\[6\] _2774_ egd_top.BitStream_buffer.buffer_index\[4\]
+ _2793_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__or4b_4
XFILLER_0_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5574_ _2278_ _2279_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4525_ _1238_ _1239_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__nand2_1
X_4456_ _0378_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__inv_2
X_4387_ _2848_ _0945_ _0946_ _0333_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__a221oi_1
X_3407_ _2933_ _2837_ vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__and2_1
X_3338_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__buf_4
X_6126_ _2693_ _2656_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__nand2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _2629_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ sky130_fd_sc_hd__inv_2
X_3269_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__buf_4
X_5008_ _0797_ _2814_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4310_ _1024_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__nand2_1
X_5290_ _0992_ _3066_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _3155_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__buf_4
X_4172_ _2953_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__buf_2
XFILLER_0_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3956_ _3001_ _3037_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5626_ _2307_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
X_3887_ _0417_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _0606_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5557_ _2261_ _2262_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__nand2_1
X_4508_ _1126_ _0956_ _0538_ _0958_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__o22ai_1
X_5488_ _0602_ _0843_ _2193_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4439_ _0816_ _3058_ _0817_ _2822_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__a221oi_1
X_6109_ _2660_ _2677_ _2661_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__nand3_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6181__50 clknet_1_1__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__inv_2
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4790_ _0816_ _3070_ _0817_ _2828_ _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__a221oi_1
X_3810_ _3039_ _3015_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__nand2_1
XANTENNA_29 _2833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3741_ net221 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_18 _1206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3672_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6460_ net202 _0293_ net43 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_5411_ egd_top.BitStream_buffer.BS_buffer\[80\] _0996_ _1000_ _0997_ _2117_ vssd1
+ vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__a221oi_1
X_6391_ net133 _0224_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_5342_ _2048_ _2049_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5273_ _0874_ _0638_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__nand2_1
X_4224_ _0397_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__clkbuf_4
X_4155_ _2976_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__clkbuf_4
X_4086_ _0802_ _3070_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4988_ _0939_ _3146_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3939_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5609_ egd_top.BitStream_buffer.buffer_index\[6\] egd_top.BitStream_buffer.buffer_index\[5\]
+ _2775_ _2793_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__or4b_4
XFILLER_0_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6233__98 clknet_1_1__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
XFILLER_0_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 la_data_in_47_32[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_4
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5960_ _2489_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__inv_2
X_4911_ _1620_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__nand2_1
X_5891_ _2467_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4842_ _1543_ _1546_ _1549_ _1553_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__and4_1
X_4773_ _0791_ _3066_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3724_ _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3655_ _0373_ egd_top.BitStream_buffer.BS_buffer\[86\] _0374_ egd_top.BitStream_buffer.BS_buffer\[87\]
+ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a22o_1
X_6443_ net185 _0276_ net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6374_ net116 _0207_ net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_3586_ _3134_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__buf_4
X_5325_ _0947_ _0371_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__nand2_1
X_6160__31 clknet_1_1__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__inv_2
X_5256_ _1953_ _1957_ _1959_ _1963_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ _0923_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _0924_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5187_ _2820_ _0954_ _2818_ _0955_ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_3_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4138_ _0444_ _2854_ _0854_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__o21ai_1
X_4069_ _0458_ _0781_ _3037_ _0782_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3440_ _2856_ _2985_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__and2_1
X_3371_ egd_top.BitStream_buffer.BS_buffer\[26\] vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__buf_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _2619_ _2565_ _2659_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__o21ai_2
X_5110_ _1781_ _1790_ _1804_ _1819_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _0865_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1751_
+ sky130_fd_sc_hd__nand2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5943_ _2481_ _2499_ _2441_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__o21ai_1
X_6282__144 clknet_1_1__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
XFILLER_0_75_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5874_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] vssd1 vssd1 vccd1 vccd1
+ _2451_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4825_ _0897_ _0495_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6212__79 clknet_1_1__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
XFILLER_0_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4756_ _0414_ _0987_ _0551_ _0989_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3707_ _2878_ _2836_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__and2_1
X_4687_ _2858_ _0657_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__nand2_1
X_6426_ net168 _0259_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_3638_ _0357_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0358_
+ sky130_fd_sc_hd__or2b_1
X_6357_ net99 _0190_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3569_ _3117_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__buf_4
X_5308_ _0602_ _3083_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__or2_1
X_5239_ _0804_ _0886_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 egd_top.BitStream_buffer.BitStream_buffer_valid_n vssd1 vssd1 vccd1 vccd1 net225
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4610_ _0925_ _0587_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5590_ _2288_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__clkbuf_1
X_4541_ _3070_ _0787_ _2922_ _0788_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4472_ _0516_ _0882_ _1183_ _1184_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3423_ _2971_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _2972_
+ sky130_fd_sc_hd__nand2_1
X_6142_ _2693_ _2656_ _2708_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__nand3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3354_ _2902_ _2852_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__and2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _2451_ _2608_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__xor2_1
X_3285_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _2834_ sky130_fd_sc_hd__inv_2
X_5024_ _0833_ _2822_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__nand2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5926_ _2500_ _2451_ _2501_ _2502_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5857_ _2435_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5788_ egd_top.BitStream_buffer.pc_reg\[5\] vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4808_ _1519_ _2912_ _1052_ _2917_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_90_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4739_ _1450_ _1451_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6409_ net151 _0242_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _0686_ _3032_ _0687_ _0688_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__o2111a_1
X_5711_ _2793_ _2779_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5642_ _2315_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5573_ net221 egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1
+ vccd1 _2279_ sky130_fd_sc_hd__nand2_1
X_4524_ _0999_ _0926_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4455_ _0495_ _2840_ _2847_ _0894_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__a221oi_1
X_4386_ _1100_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3406_ _2944_ _2945_ _2948_ _2950_ _2954_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__o2111a_1
X_6125_ _2689_ _2674_ _2512_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__o21ai_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _2885_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__buf_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _2615_ _2560_ _2488_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__or3_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _2821_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__clkbuf_1
X_5007_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__inv_2
X_3199_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5909_ _2458_ _2475_ _2473_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6333__23 clknet_1_0__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__inv_2
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4240_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__inv_2
X_4171_ _3139_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ _2999_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _0673_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6167__37 clknet_1_1__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__inv_2
X_5625_ net15 _3017_ _2299_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__mux2_1
X_3886_ _0603_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5556_ _0949_ _0709_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__nand2_1
X_4507_ _1210_ _1213_ _1217_ _1221_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__and4_2
X_5487_ _0844_ _3066_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4438_ _1151_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__nand2_1
X_4369_ _2944_ _3084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__or2_1
X_6108_ _2675_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__inv_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _2496_ _2607_ _2610_ _2489_ _2613_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__o221a_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ _3074_ _0453_ _0457_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__a31o_1
XANTENNA_19 _1495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3671_ _2902_ _2937_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__and2_1
X_5410_ _2115_ _2116_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__nand2_1
X_6390_ net132 _0223_ net50 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5341_ _2881_ _0456_ _2790_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__o21a_1
X_5272_ _2951_ _0863_ _0864_ _0385_ _1979_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__a221oi_2
X_4223_ _0939_ _0341_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__nand2_1
X_4154_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4085_ _3057_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4987_ _0894_ _0945_ _0946_ egd_top.BitStream_buffer.BS_buffer\[46\] _1697_ vssd1
+ vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_73_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3938_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__clkbuf_8
X_3869_ _0373_ egd_top.BitStream_buffer.BS_buffer\[87\] _0374_ _0587_ vssd1 vssd1
+ vccd1 vccd1 _0588_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5608_ _2297_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
X_5539_ _3086_ _2957_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 la_data_in_49_48[0] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4910_ _0835_ _1011_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__nand2_1
X_5890_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _2952_ _3077_ _1550_ _1551_ _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4772_ _2874_ _0781_ _3153_ _0782_ _1483_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3723_ egd_top.BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__buf_4
X_6442_ net184 _0275_ net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3654_ _2893_ _2852_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6373_ net115 _0206_ net41 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3585_ _2845_ _2910_ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5324_ _0937_ _0553_ _2859_ _0938_ _2031_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5255_ _0607_ _0831_ _0832_ _0625_ _1962_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__a221oi_1
X_4206_ _0357_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5186_ _3067_ _0956_ _1372_ _0958_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_3_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4137_ _2858_ _2848_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ egd_top.BitStream_buffer.BS_buffer\[126\] _0783_ _0784_ _2828_ vssd1 vssd1
+ vccd1 vccd1 _0785_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3370_ _2856_ _2915_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__and2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _1741_ _1744_ _1747_ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5942_ _2517_ _2518_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5873_ _2448_ _2449_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4824_ _0895_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _1536_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4755_ _1466_ _1467_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3706_ _0418_ _0421_ _0423_ _0425_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4686_ _3010_ _0848_ _3017_ _0849_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6425_ net167 _0258_ net39 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_3637_ _2870_ _2852_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6356_ net98 _0189_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3568_ _2933_ _2937_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5307_ _0984_ _3079_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__or2_1
X_3499_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__buf_4
X_5238_ _0802_ _2812_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__nand2_1
X_5169_ _0889_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _1878_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6266__129 clknet_1_0__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__2731_ clknet_0__2731_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2731_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4540_ _3154_ _0790_ _1253_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4471_ _1185_ _0889_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3422_ _2902_ _2837_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__and2_1
X_6141_ _2704_ _2505_ _2562_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__nand3_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _2898_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__and3_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _2832_ _2764_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__nor2_4
X_6072_ _2454_ _2640_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__nor2_1
X_5023_ _0824_ _2907_ _0825_ _3127_ _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__a221oi_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1 vccd1 vccd1
+ _2502_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5856_ net8 _2904_ _2419_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4807_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5787_ _2393_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
X_4738_ _0949_ _0366_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4669_ _2800_ _0810_ _2990_ _0809_ _1381_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6408_ net150 _0241_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6339_ net81 _0172_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[91\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188__57 clknet_1_0__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__inv_2
XFILLER_0_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3971_ _3039_ _3017_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5710_ _2351_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
X_5641_ net1 _3090_ _2298_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5572_ _2276_ _2277_ vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4523_ _0428_ _0657_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4454_ _0772_ _2854_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4385_ _0949_ _3142_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3405_ _2952_ _2953_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__or2_1
X_6124_ _2680_ _2691_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__nand2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _2884_ _2865_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__and2_1
X_6055_ _2628_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ sky130_fd_sc_hd__inv_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _2802_ _0787_ _3090_ _0788_ _1715_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__a221oi_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ net11 _2820_ _2797_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__mux2_1
X_6249__113 clknet_1_1__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
X_3198_ _2766_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__buf_6
XFILLER_0_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5908_ _2484_ _2471_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5839_ _2426_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4170_ _0885_ _0886_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3954_ _2997_ _2816_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3885_ _0411_ _0414_ _0413_ _2887_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a22o_1
X_5624_ _2306_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__clkbuf_1
X_5555_ _0947_ _3105_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5486_ _2181_ _2185_ _2187_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__and4_1
X_4506_ _0464_ _0945_ _0946_ _3143_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__a221oi_1
X_4437_ _0820_ _2814_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6107_ _2662_ _2675_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__nand2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _0650_ _3080_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_1
X_4299_ egd_top.BitStream_buffer.BS_buffer\[127\] _0783_ _0784_ _0458_ vssd1 vssd1
+ vccd1 vccd1 _1015_ sky130_fd_sc_hd__a22o_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__inv_2
X_6038_ _2611_ _2612_ _2500_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__o21ai_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3670_ _0388_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5340_ _1994_ _0903_ _2047_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__nand3_1
X_5271_ _1977_ _1978_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__nand2_1
X_4222_ _0394_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__clkbuf_4
X_4153_ _3119_ _0863_ _0864_ _0346_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__a221oi_2
X_4084_ _3056_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4986_ _1695_ _1696_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3937_ _0650_ _2945_ _0651_ _0652_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__o2111a_1
X_3868_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5607_ net1 _0414_ _2280_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__mux2_1
X_3799_ _3014_ _3017_ _3016_ _0402_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a22o_1
X_5538_ _0984_ _3083_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5469_ _0804_ _0469_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__nand2_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 la_data_in_49_48[1] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4840_ _3087_ _0392_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4771_ egd_top.BitStream_buffer.BS_buffer\[3\] _0783_ _0784_ _0886_ vssd1 vssd1 vccd1
+ vccd1 _1483_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3722_ _0439_ egd_top.BitStream_buffer.BS_buffer\[90\] _0441_ egd_top.BitStream_buffer.BS_buffer\[91\]
+ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6441_ net183 _0274_ net42 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3653_ _2899_ _2852_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__and2_1
X_6372_ net114 _0205_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_3584_ _3132_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__inv_2
X_5323_ _2029_ _2030_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__nand2_1
X_5254_ _1960_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__nand2_1
X_5185_ _1883_ _1886_ _1889_ _1893_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__and4_1
X_4205_ _0363_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _0414_ _0848_ _3010_ _0849_ _0852_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4067_ _3044_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4969_ _0990_ _3048_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5941_ _2505_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1
+ vccd1 _2518_ sky130_fd_sc_hd__nand2_1
X_6243__108 clknet_1_1__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5872_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] vssd1 vssd1 vccd1 vccd1
+ _2449_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4823_ _0602_ _0882_ _1531_ _1532_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4754_ _0992_ _3030_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _0424_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _0425_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4685_ _0544_ _0850_ _1397_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__o21ai_1
X_3636_ _3150_ _0332_ _0345_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__and4_1
X_6424_ net166 _0257_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_3567_ _3114_ _3115_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__nand2_1
X_6355_ net97 _0188_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5306_ _3143_ _3095_ _3103_ egd_top.BitStream_buffer.BS_buffer\[83\] _2013_ vssd1
+ vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__a221oi_2
X_5237_ _2824_ _2996_ _2927_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__a31oi_1
X_3498_ _3046_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5168_ _0885_ _2881_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__nand2_1
X_4119_ _0835_ _2824_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__nand2_1
X_5099_ _0949_ _0371_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__2730_ clknet_0__2730_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2730_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6202__70 clknet_1_1__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__inv_2
XFILLER_0_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4470_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3421_ _2969_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _2970_
+ sky130_fd_sc_hd__nand2_1
X_6140_ _2694_ _2706_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__nand2_1
X_3352_ _2900_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _2901_
+ sky130_fd_sc_hd__nand2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _2831_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__nand2_4
XFILLER_0_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6071_ _2640_ _2454_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _0983_ _0826_ _2981_ _0827_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__o22ai_1
X_5924_ _2477_ _2491_ _2466_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__nor3_1
X_5855_ _2434_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _1000_ _2840_ _2847_ _0926_ _1517_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__a221oi_1
X_5786_ net1 _0330_ _2376_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4737_ _0947_ _3139_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4668_ _1052_ _0811_ _1380_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__o21ai_1
X_3619_ _0334_ _0335_ _0337_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__o22ai_1
X_6407_ net149 _0240_ net49 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_4599_ _2952_ _3110_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__o21ai_1
X_6338_ net80 _0171_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[92\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6272__134 clknet_1_1__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _3036_ _2990_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _2314_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5571_ _0412_ _0456_ _2789_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__o21a_1
X_4522_ _2943_ _0987_ _0841_ _0989_ _1236_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4453_ _2858_ _2959_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__nand2_1
X_3404_ _2845_ _2769_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__nand2_1
X_4384_ _0947_ _2951_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nand2_1
X_6123_ _2690_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__inv_2
X_3335_ _2883_ _2875_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__nor2_8
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _2615_ _2560_ _2478_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__or3_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__buf_6
X_5005_ _3064_ _0790_ _1714_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__o21ai_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3197_ _2765_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5907_ _2483_ _2443_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] egd_top.BitStream_buffer.BitStream_buffer_output\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5838_ net2 _0926_ _2420_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5769_ _2384_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_6193__61 clknet_1_0__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__inv_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6295__156 clknet_1_1__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__inv_2
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3953_ _3091_ _2982_ _0668_ _0669_ _0670_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__o2111a_1
X_3884_ _0601_ _0405_ _0602_ _0409_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5623_ net16 _3015_ _2299_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5554_ _0937_ _2859_ _0463_ _0938_ _2259_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__a221oi_1
X_6324__14 clknet_1_1__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__inv_2
X_5485_ _0477_ _0831_ _0832_ _1011_ _2190_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__a221oi_1
X_4505_ _1218_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__nand2_1
X_4436_ _0818_ _2820_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4367_ _3124_ _3096_ _3104_ _2830_ _1082_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__a221oi_2
X_6106_ _2674_ _2512_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _2866_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__clkbuf_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _1013_ _1014_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__nand2_1
X_3249_ net2 _2808_ _2798_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__mux2_1
X_6037_ _2453_ _2578_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6303__163 clknet_1_1__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__inv_2
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6278__140 clknet_1_0__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
X_6172__42 clknet_1_0__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__inv_2
X_5270_ _0867_ _0389_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4221_ _0391_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__buf_4
X_4152_ _0866_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nand2_1
X_4083_ _3055_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4985_ _0949_ _2957_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3936_ _0653_ _2953_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__or2_1
X_3867_ _0435_ _0368_ _0370_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1
+ vccd1 vccd1 _0586_ sky130_fd_sc_hd__a22o_1
X_5606_ _2296_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__clkbuf_1
X_3798_ _0516_ _3009_ _0407_ _3012_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5537_ _0601_ _3079_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__or2_1
X_5468_ _0802_ _2816_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5399_ _0756_ _0882_ _2103_ _2104_ _2105_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__o2111a_1
X_4419_ _1133_ _1134_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__nand2_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 la_data_in_65 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6209__76 clknet_1_1__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4770_ _1481_ _1482_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__nand2_1
X_3721_ _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__clkbuf_4
X_6440_ net182 _0273_ net41 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3652_ _0366_ _0368_ _0370_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a22o_1
X_6371_ net113 _0204_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_3583_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__buf_4
XFILLER_0_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5322_ _0941_ _2848_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5253_ _0835_ _0469_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__nand2_1
X_5184_ _0888_ _3077_ _1890_ _1891_ _1892_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__o2111a_1
X_4204_ _0361_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__clkbuf_4
X_4135_ _0474_ _0850_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4066_ _3043_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4968_ _0981_ _3017_ _0982_ _0402_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4899_ _1599_ _1602_ _1605_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3919_ _2900_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0637_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6316__7 clknet_1_1__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__inv_2
XFILLER_0_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5940_ _2516_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1
+ vccd1 _2517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5871_ _2446_ _2447_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__nand2_1
X_4822_ _1533_ _0889_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__or2_1
X_4753_ _0990_ _2987_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3704_ _2884_ _2984_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6423_ net165 _0256_ net41 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_4684_ _2867_ _2907_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3635_ _0351_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__nor2_1
X_6354_ net96 _0187_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3566_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__buf_4
X_5305_ _0337_ _3092_ _2012_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__o21ai_1
X_3497_ _2870_ _2984_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__nand2_1
X_5236_ _1372_ _0796_ _1943_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5167_ _0883_ _2943_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4118_ _3026_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__clkbuf_4
X_5098_ _0947_ _0435_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__nand2_1
X_4049_ _0430_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _0767_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3420_ _2933_ _2852_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3351_ _2899_ _2872_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ egd_top.BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__inv_2
X_6070_ _2542_ _2531_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__nand2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _0816_ _2791_ _0817_ _0625_ _1730_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__a221oi_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5923_ _2477_ _2499_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5854_ net9 _0607_ _2419_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4805_ _3031_ _2854_ _1516_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5785_ _2392_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
X_4736_ _0937_ _0435_ _0371_ _0938_ _1448_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4667_ _0812_ _2863_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__nand2_1
X_6406_ net148 _0239_ net52 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_3618_ _2833_ _2910_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6337_ net79 _0170_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[93\]
+ sky130_fd_sc_hd__dfrtp_2
X_4598_ _3118_ _3115_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__nand2_1
X_3549_ _3096_ _3097_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__nand2_1
X_5219_ _0937_ _3105_ _0709_ _0938_ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5570_ _2222_ _0903_ _2275_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__nand3_2
XFILLER_0_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4521_ _1234_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4452_ _3007_ _0848_ _3040_ _0849_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__a221oi_1
X_3403_ _2951_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4383_ _0937_ _3139_ _0366_ _0938_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6122_ _2689_ _2512_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__nand2_1
X_3334_ _2831_ _2868_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__nand2_8
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _2625_ _2627_ vssd1 vssd1 vccd1 vccd1 egd_top.exp_golomb_decoding.te_range\[2\]
+ sky130_fd_sc_hd__nor2_1
X_3265_ _2819_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _0791_ _3070_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__nand2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _2764_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] egd_top.BitStream_buffer.BitStream_buffer_output\[2\]
+ _2441_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__o21a_1
X_5837_ _2425_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5768_ net16 _3002_ _2377_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__mux2_1
X_4719_ _1287_ _3093_ _1431_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5699_ net12 _3115_ _2335_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3952_ _2992_ _0406_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3883_ _3040_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5622_ _2305_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__clkbuf_1
X_5553_ _2257_ _2258_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__nand2_1
X_4504_ _0949_ _3139_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5484_ _2188_ _2189_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4435_ _3037_ _0809_ _0330_ _0810_ _1149_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4366_ _0859_ _3093_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o21ai_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _2671_ _2673_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__nand2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _2864_ _2865_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__and2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1
+ vccd1 vccd1 _1014_ sky130_fd_sc_hd__nand2_1
X_3248_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__buf_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _2455_ _2532_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__nor2_1
X_3179_ net30 net29 vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6158__29 clknet_1_0__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__inv_2
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4220_ _0388_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _0867_ _3112_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__nand2_1
X_4082_ _0795_ _3065_ _0723_ _0796_ _0798_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__o221a_1
X_4984_ _0947_ _0366_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__nand2_1
X_3935_ _3142_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5605_ net8 _0412_ _2280_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__mux2_1
X_3866_ _0580_ _0581_ _0582_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3797_ _2993_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__inv_2
X_5536_ _3146_ _3095_ _3103_ egd_top.BitStream_buffer.BS_buffer\[85\] _2241_ vssd1
+ vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__a221oi_2
X_5467_ _2828_ _2996_ _2927_ _2172_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__a31oi_1
X_4418_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] vssd1 vssd1
+ vccd1 vccd1 _1134_ sky130_fd_sc_hd__nand2_1
X_5398_ _0889_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _2105_
+ sky130_fd_sc_hd__or2b_1
X_4349_ _0885_ _2874_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nand2_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6019_ _2593_ _2590_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3720_ _2833_ _2851_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__clkbuf_8
X_6370_ net112 _0203_ net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3582_ _3130_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__clkbuf_4
X_5321_ _0939_ _2931_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__nand2_1
X_5252_ _0833_ _2826_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5183_ _3087_ _0398_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__nand2_1
X_4203_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4134_ _2867_ _2913_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4065_ _3047_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _0480_ _0405_ _2981_ _0409_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__o22ai_1
X_4898_ _2802_ _0800_ _0801_ _2824_ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__a221oi_1
X_3918_ _2896_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _0636_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3849_ _0444_ _3152_ _0567_ _3155_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5519_ _0990_ _2990_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6499_ net73 _0325_ net35 vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2729_ clknet_0__2729_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2729_
+ sky130_fd_sc_hd__clkbuf_16
X_5870_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] vssd1 vssd1 vccd1 vccd1
+ _2447_ sky130_fd_sc_hd__inv_2
X_4821_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4752_ _0981_ _3040_ _0982_ _3015_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__a221oi_1
X_3703_ _0422_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0423_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4683_ _3101_ _0840_ _2943_ _0842_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3634_ _0352_ egd_top.BitStream_buffer.BS_buffer\[126\] _0353_ egd_top.BitStream_buffer.BS_buffer\[127\]
+ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__a22o_1
X_6422_ net164 _0255_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3565_ _2856_ _2937_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6353_ net95 _0186_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_5304_ _3099_ _3015_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__nand2_1
X_3496_ egd_top.BitStream_buffer.BS_buffer\[123\] _3043_ _3044_ egd_top.BitStream_buffer.BS_buffer\[124\]
+ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__a22o_1
X_5235_ _0797_ _2818_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _0892_ _2959_ _0893_ _0583_ _1874_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__a221oi_1
X_4117_ _0833_ _2808_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__nand2_1
X_5097_ _2987_ _0922_ _0607_ _0921_ _1806_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4048_ _0428_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _0766_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5999_ _2570_ _2574_ _2509_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__nand3_1
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3350_ _2898_ egd_top.BitStream_buffer.pc\[2\] _2868_ vssd1 vssd1 vccd1 vccd1 _2899_
+ sky130_fd_sc_hd__and3_4
XFILLER_0_29_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _1728_ _1729_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__nand2_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__buf_4
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ _2464_ _2491_ _2465_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__nand3_4
XFILLER_0_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5853_ _2433_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5784_ net8 _3070_ _2376_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__mux2_1
X_4804_ _2858_ _0894_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__nand2_1
X_4735_ _1446_ _1447_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4666_ _1368_ _1371_ _1374_ _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__and4_1
X_6405_ net147 _0238_ net52 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_3617_ _0336_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
X_4597_ _0343_ _3126_ _2974_ _3123_ _1310_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__a221oi_1
X_6336_ net78 _0169_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[94\]
+ sky130_fd_sc_hd__dfrtp_4
X_3548_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3479_ _3021_ _3023_ _3025_ _3027_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__and4_1
X_5218_ _1925_ _1926_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__nand2_1
X_5149_ _2858_ _0926_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4520_ _0992_ _3048_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4451_ _0546_ _0850_ _1165_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__o21ai_1
X_3402_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__buf_4
X_6121_ _2681_ _2688_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__nor2_1
X_4382_ _1096_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nand2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _2880_ _2881_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__nand2_1
X_6052_ _2626_ _2557_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__nand2_1
X_3264_ net12 _2818_ _2798_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__mux2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _0988_ _0781_ _0330_ _0782_ _1712_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__a221oi_1
X_3195_ egd_top.BitStream_buffer.pc\[0\] egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1
+ vccd1 vccd1 _2764_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5905_ _2481_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5836_ net3 _0830_ _2420_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5767_ _2383_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
X_5698_ _2345_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
X_4718_ _3100_ _3007_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4649_ _1309_ _0903_ _1362_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _2989_ _3066_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3882_ _2863_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5621_ net2 _3040_ _2299_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5552_ _0941_ _2959_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4503_ _0947_ _0392_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5483_ _0835_ _1116_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4434_ _0641_ _0811_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__o21ai_1
X_4365_ _3100_ _0412_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6104_ _2532_ _2608_ _2533_ _2672_ _2489_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__a311o_1
X_3316_ _2768_ _2835_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _2865_
+ sky130_fd_sc_hd__and3_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _2608_ _2609_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__nor2_1
X_4296_ _1010_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nand2_1
X_3247_ _2807_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__clkbuf_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _2744_ net28 vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__nand2_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5819_ net35 egd_top.BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6239__104 clknet_1_0__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XFILLER_0_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4150_ _2938_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__clkbuf_4
X_4081_ _0797_ _2800_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6285__146 clknet_1_1__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__inv_2
X_4983_ _0443_ _0922_ _0420_ _0921_ _1693_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__a221oi_1
X_3934_ _2949_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _0652_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3865_ _0363_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5604_ _2295_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
X_3796_ _0511_ _0512_ _0513_ _0514_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5535_ _3133_ _3092_ _2240_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__o21ai_1
X_5466_ _1603_ _0796_ _2171_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ _1131_ _1132_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5397_ _0885_ _0412_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__nand2_1
X_4348_ _0883_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _1064_
+ sky130_fd_sc_hd__nand2_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4279_ _0434_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__clkbuf_4
X_6018_ _2552_ _2589_ _2514_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3581_ _2964_ _2937_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__nand2_1
X_5320_ _3048_ _0922_ _0477_ _0921_ _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__a221oi_1
X_5251_ _0824_ _3124_ _0825_ _0395_ _1958_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_11_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4202_ _0906_ _0911_ _0914_ _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__and4_1
X_5182_ _0407_ _3084_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4133_ _0629_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__clkbuf_4
X_4064_ _3050_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ _1670_ _1672_ _1674_ _1676_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__and4_1
X_4897_ _1606_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__nand2_1
X_3917_ _2848_ _2839_ _2846_ _2959_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3848_ _3070_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3779_ _0496_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5518_ _0981_ _2913_ _0982_ _2980_ _2223_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__a221oi_1
X_6498_ net72 egd_top.BitStream_buffer.pc\[6\] net35 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_5449_ _0653_ _0969_ _0904_ _0971_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6214__81 clknet_1_1__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2728_ clknet_0__2728_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2728_
+ sky130_fd_sc_hd__clkbuf_16
X_4820_ _0885_ _0841_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4751_ _3091_ _0405_ _0983_ _0409_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__o22ai_1
X_3702_ _2964_ _2871_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4682_ _0489_ _0843_ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__o21ai_1
X_3633_ _2767_ _2996_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__and2_1
X_6421_ net163 _0254_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3564_ _3111_ _3112_ vssd1 vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__nand2_1
X_6352_ net94 _0185_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6283_ clknet_1_0__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__buf_1
X_5303_ _3142_ _0907_ _0656_ _0908_ _2010_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__a221oi_1
X_3495_ _2878_ _2961_ vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__and2_1
X_5234_ _2806_ _0787_ _3127_ _0788_ _1941_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__a221oi_1
X_5165_ _1872_ _1873_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _3024_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5096_ _2849_ _0923_ _1805_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o21ai_1
X_4047_ _0761_ _0762_ _0763_ _0764_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5998_ _2508_ _2522_ _2573_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__nand3_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4949_ _0389_ _0907_ _0435_ _0908_ _1659_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3280_ _2829_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__clkbuf_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _2490_ _2497_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5852_ net10 _0420_ _2419_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5783_ _2391_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4803_ _0406_ _0848_ _0402_ _0849_ _1514_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__a221oi_1
X_4734_ _0941_ _0553_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4665_ _2791_ _0800_ _0801_ _2820_ _1377_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6404_ net146 _0237_ net52 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_4596_ _0492_ _3131_ _0574_ _3135_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__o22ai_1
X_3616_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6335_ net77 _0168_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_3547_ _3095_ vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3478_ _3026_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _3027_
+ sky130_fd_sc_hd__nand2_1
X_5217_ _0941_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _1926_
+ sky130_fd_sc_hd__nand2_1
X_5148_ _3017_ _0848_ _2922_ _0849_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__a221oi_1
X_5079_ _0974_ _2939_ _0975_ _2926_ _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_66_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4450_ _2867_ _3097_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4381_ _0941_ _0371_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__nand2_1
X_3401_ _2949_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _2950_
+ sky130_fd_sc_hd__nand2_1
X_6120_ _2686_ _2687_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__nand2_1
X_3332_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__clkbuf_8
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _2622_ _2624_ _2623_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__nand3_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__clkbuf_8
X_3194_ _2763_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[0\] sky130_fd_sc_hd__clkinv_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ egd_top.BitStream_buffer.BS_buffer\[5\] _0783_ _0784_ _0469_ vssd1 vssd1 vccd1
+ vccd1 _1712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5904_ _2479_ _2480_ vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__nand2_4
X_5835_ _2424_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5766_ net2 _3048_ _2377_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__mux2_1
X_5697_ net13 egd_top.BitStream_buffer.BS_buffer\[57\] _2335_ vssd1 vssd1 vccd1 vccd1
+ _2345_ sky130_fd_sc_hd__mux2_1
X_4717_ _3115_ _0907_ _0398_ _0908_ _1429_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4648_ _1322_ _1338_ _1347_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__and4_1
X_4579_ _1291_ _1292_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6184__53 clknet_1_1__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__inv_2
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3950_ _2986_ _3048_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__nand2_1
X_3881_ _0585_ _0589_ _0594_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__and4_2
XFILLER_0_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5620_ _2304_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__clkbuf_1
X_5551_ _0939_ _2926_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__nand2_1
X_4502_ _0937_ _0398_ _0435_ _0938_ _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__a221oi_1
X_5482_ _0833_ _0458_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4433_ _0812_ _3017_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4364_ egd_top.BitStream_buffer.BS_buffer\[55\] _0907_ _0392_ _0908_ _1079_ vssd1
+ vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__a221oi_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _2832_ _2842_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__nor2_4
X_6103_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] _2608_ vssd1 vssd1
+ vccd1 vccd1 _2672_ sky130_fd_sc_hd__nor2_1
X_4295_ _1011_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__o21a_1
X_3246_ net3 _2806_ _2798_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__mux2_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _2449_ _2469_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__nor2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3177_ _2742_ _2743_ _2745_ _2746_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6262__125 clknet_1_1__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5818_ _2415_ _2398_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[2\] sky130_fd_sc_hd__xnor2_4
X_5749_ _2795_ _2372_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ _3069_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4982_ _0620_ _0923_ _1692_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3933_ _2947_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0651_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3864_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5603_ net9 _2943_ _2280_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__mux2_1
X_3795_ _3004_ _2806_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5534_ _3099_ _0402_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__nand2_1
X_5465_ _0797_ _2822_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__nand2_1
X_6163__34 clknet_1_1__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__inv_2
XFILLER_0_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4416_ _0886_ _0457_ _2790_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__o21a_1
X_5396_ _0883_ _0414_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__nand2_1
X_4347_ _0420_ _0872_ _0894_ _0873_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__a221oi_1
X_4278_ _0551_ _0987_ _0988_ _0989_ _0994_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__a221oi_2
X_3229_ net224 egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1
+ _2794_ sky130_fd_sc_hd__nand2_1
X_6017_ _2552_ _2565_ _2592_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__o21ai_2
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3580_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5250_ _2981_ _0826_ _3091_ _0827_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__o22ai_1
X_4201_ _3129_ _3077_ _0915_ _0916_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__o2111a_1
X_5181_ _0757_ _3080_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _2886_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__clkbuf_4
X_4063_ _0779_ _0780_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4965_ _0974_ _2931_ _0975_ _2939_ _1675_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3916_ _3151_ _2853_ _0633_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4896_ _0804_ _0625_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__nand2_1
X_3847_ _0398_ _3141_ _2771_ _3139_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _2965_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _0497_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5517_ _1287_ _0404_ _0641_ _0408_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__o22ai_1
X_6497_ net71 egd_top.BitStream_buffer.pc\[5\] net36 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5448_ _2848_ _0961_ _0962_ _0463_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__a221oi_1
X_5379_ _3067_ _2853_ _2085_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__o21ai_1
X_6268__131 clknet_1_0__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_0_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2727_ clknet_0__2727_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2727_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4750_ _1456_ _1458_ _1460_ _1462_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3701_ _0419_ _0420_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_1
X_4681_ _0844_ _3048_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__nand2_1
X_3632_ _2902_ _2996_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__and2_1
X_6420_ net162 _0253_ net40 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6351_ net93 _0184_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3563_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__buf_4
X_5302_ _1301_ _3109_ _2009_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__o21ai_1
X_3494_ _2833_ _2961_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__and2_1
X_5233_ _0698_ _0790_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5164_ _0897_ _1000_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__nand2_1
X_4115_ _3020_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__clkbuf_4
X_5095_ _0925_ _0420_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__nand2_1
X_4046_ _0424_ _0443_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5997_ _2571_ _2572_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4948_ _0888_ _3110_ _1658_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__o21ai_1
X_4879_ _1589_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5920_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _2494_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ _2496_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__o22ai_1
X_5851_ _2432_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5782_ net9 _3153_ _2376_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__mux2_1
X_4802_ _2944_ _0850_ _1513_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__o21ai_1
X_4733_ _0939_ _3143_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6403_ net145 _0236_ net52 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[53\]
+ sky130_fd_sc_hd__dfrtp_4
X_4664_ _1375_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3615_ _2864_ _2910_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4595_ _1263_ _1277_ _1290_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3546_ _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__clkbuf_2
X_5216_ _0939_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1925_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3477_ _2856_ _2961_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__and2_1
X_5147_ _0881_ _0850_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__o21ai_1
X_5078_ _0574_ _0976_ _3075_ _0977_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__o22ai_1
X_4029_ _0382_ _0385_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2729_ _2729_ vssd1 vssd1 vccd1 vccd1 clknet_0__2729_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4380_ _0939_ _0343_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__nand2_1
X_3400_ _2927_ _2872_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__and2_1
X_3331_ _2879_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__buf_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _2622_ _2623_ _2624_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__a21oi_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _2817_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__clkbuf_1
X_3193_ _2761_ _2762_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__nand2_4
X_5001_ _1710_ _1711_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__nand2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5903_ _2471_ _2474_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__nand2_2
X_5834_ net4 _1000_ _2420_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5765_ _2382_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5696_ _2344_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4716_ _0492_ _3110_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__o21ai_1
X_4647_ _1349_ _1353_ _1357_ _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4578_ _0867_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _1292_
+ sky130_fd_sc_hd__nand2_1
X_3529_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__inv_2
X_6179_ clknet_1_0__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__buf_1
XFILLER_0_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3880_ _0595_ _0596_ _0597_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5550_ _0610_ _0921_ _3030_ _0922_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5481_ _0824_ _2935_ _0825_ _0378_ _2186_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__a221oi_1
X_4501_ _1214_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4432_ _1136_ _1139_ _1142_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4363_ _0904_ _3110_ _1078_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__o21ai_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6102_ _2669_ _2670_ _2509_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__nand3_1
X_3314_ egd_top.BitStream_buffer.BS_buffer\[25\] vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__buf_4
X_4294_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__clkbuf_8
X_3245_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__buf_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _2468_ _2543_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__nor2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _2743_ net29 vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5817_ _2399_ _2400_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5748_ _2794_ _2774_ vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__nand2_1
X_5679_ net7 _2939_ _2335_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4981_ _0925_ _0871_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _0414_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__inv_2
X_3863_ _0361_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0582_
+ sky130_fd_sc_hd__nand2_1
X_5602_ _2294_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__clkbuf_1
X_3794_ _3001_ _3030_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5533_ _0398_ _0907_ _0553_ _0908_ _2238_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _2810_ _0787_ _0395_ _0788_ _2169_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5395_ _0892_ _0657_ _0893_ _0420_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__a221oi_1
X_4415_ _1074_ _0903_ _1130_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__nand3_1
X_4346_ _1060_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nand2_1
X_4277_ _0991_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nand2_1
X_6016_ _2562_ _2551_ _2588_ _2591_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__a31o_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _2745_ _2749_ _2737_ net223 vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__a22o_2
X_3159_ net32 net31 vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6291__152 clknet_1_0__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__inv_2
X_4200_ _3087_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0917_
+ sky130_fd_sc_hd__nand2_1
X_5180_ _0333_ _3096_ _3104_ _0894_ _1888_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__a221oi_1
X_4131_ _2880_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4062_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1
+ vccd1 vccd1 _0780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4964_ _0347_ _0976_ _0730_ _0977_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3915_ _2857_ _0463_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4895_ _0802_ _2806_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3846_ _0337_ _3145_ _3133_ _3148_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3777_ _2962_ _2818_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__nand2_1
X_6496_ net70 egd_top.BitStream_buffer.pc\[4\] net36 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5516_ _2178_ _2192_ _2204_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5447_ _3108_ _0963_ _0561_ _0964_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__o22ai_1
X_5378_ _2857_ _0875_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__nand2_1
X_4329_ _0988_ _0840_ _3101_ _0842_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__2726_ clknet_0__2726_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2726_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3700_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__buf_6
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4680_ _1382_ _1386_ _1388_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__and4_1
X_3631_ _0347_ _0348_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__o22ai_1
X_6220__86 clknet_1_0__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
X_6350_ net92 _0183_ net47 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[80\]
+ sky130_fd_sc_hd__dfrtp_2
X_3562_ _2895_ _2769_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__and2_2
XFILLER_0_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5301_ _3117_ _3139_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3493_ _3031_ _3032_ _3035_ _3038_ _3041_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__o2111a_1
X_5232_ _0791_ _2791_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__nand2_1
X_5163_ _0895_ _0886_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__nand2_1
X_4114_ _3022_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__clkbuf_4
X_5094_ _1792_ _1796_ _1800_ _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__and4_1
X_4045_ _0422_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0763_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _2515_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] _2482_ vssd1
+ vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4947_ _3118_ _2951_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__nand2_1
X_4878_ _0933_ _2904_ _0934_ _0477_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6298__158 clknet_1_0__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__inv_2
X_3829_ _3087_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _0548_
+ sky130_fd_sc_hd__nand2_1
X_6479_ net53 _0312_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5850_ net11 _0871_ _2420_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5781_ _2390_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
X_4801_ _2867_ _3127_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__nand2_1
X_4732_ _1443_ _1444_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4663_ _0804_ _2828_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3614_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__inv_2
X_6402_ net144 _0235_ net52 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[54\]
+ sky130_fd_sc_hd__dfrtp_4
X_4594_ _1294_ _1298_ _1303_ _1307_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3545_ _2902_ _2865_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__and2_1
X_3476_ _3024_ _2802_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5215_ _0830_ _0945_ _0946_ _2939_ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5146_ _2867_ _2935_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__nand2_1
X_5077_ _0967_ _1116_ _0968_ _0841_ _1786_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__a221oi_1
X_4028_ _0380_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _0746_
+ sky130_fd_sc_hd__nand2_1
X_5979_ net17 net18 vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2728_ _2728_ vssd1 vssd1 vccd1 vccd1 clknet_0__2728_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3330_ _2878_ _2871_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ net13 _2816_ _2798_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__mux2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _0461_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1
+ vccd1 _1711_ sky130_fd_sc_hd__nand2_1
X_3192_ _2760_ egd_top.BitStream_buffer.pc_reg\[0\] vssd1 vssd1 vccd1 vccd1 _2762_
+ sky130_fd_sc_hd__nand2_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5902_ _2478_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__inv_2
X_5833_ _2423_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5764_ net3 _3034_ _2377_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5695_ net14 egd_top.BitStream_buffer.BS_buffer\[56\] _2335_ vssd1 vssd1 vccd1 vccd1
+ _2344_ sky130_fd_sc_hd__mux2_1
X_4715_ _3118_ _0385_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4646_ _1358_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4577_ _0865_ _3143_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3528_ _3076_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__clkbuf_4
X_3459_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__inv_2
X_5129_ _0812_ _2980_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5480_ _3091_ _0826_ _0480_ _0827_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__o22ai_1
X_4500_ _0941_ _0656_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4431_ _3070_ _0800_ _0801_ _2816_ _1145_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__a221oi_1
XANTENNA_1 _0395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4362_ _3118_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _1078_
+ sky130_fd_sc_hd__nand2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6101_ _2637_ _2635_ _2667_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3313_ _2830_ _2840_ _2847_ _2848_ _2861_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__a221oi_2
X_4293_ _0902_ _0903_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__nand3_1
X_3244_ _2805_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__clkbuf_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _2543_ _2534_ _2606_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__o21ai_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _2742_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__nand2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5816_ _2414_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5747_ _2371_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _2334_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4629_ _3129_ _0969_ _0730_ _0971_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4980_ _1679_ _1683_ _1687_ _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__and4_1
X_3931_ _3112_ _2929_ _2930_ _2926_ _0648_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3862_ _0359_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _0581_
+ sky130_fd_sc_hd__nand2_1
X_5601_ net10 _2881_ _2280_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__mux2_1
X_3793_ _2999_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _0512_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5532_ _1533_ _3109_ _2237_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5463_ _1021_ _0790_ _2168_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5394_ _2099_ _2100_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4414_ _1088_ _1104_ _1113_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6320__11 clknet_1_0__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
X_4345_ _0877_ _3146_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__nand2_1
X_4276_ _0992_ _2987_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__nand2_1
X_6015_ _2590_ _2554_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__nand2_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _2735_ _2734_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__nand2_1
X_3158_ net33 vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6226__92 clknet_1_1__leaf__2723_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
XFILLER_0_49_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6154__25 clknet_1_0__leaf__2718_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__inv_2
XFILLER_0_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _0469_ _0840_ _0841_ _0842_ _0846_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__a221oi_1
X_4061_ _0702_ _0776_ _0457_ _0778_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4963_ _0967_ _0988_ _0968_ _1116_ _1673_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3914_ _0412_ _2880_ _2993_ _2886_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__a221oi_1
X_4894_ _1603_ _3065_ _1021_ _0796_ _1604_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3845_ _0549_ _0555_ _0559_ _0563_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__and4_1
X_3776_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6495_ net69 egd_top.BitStream_buffer.pc\[3\] net36 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5515_ _2208_ _2212_ _2216_ _2220_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ _2824_ _0954_ _2822_ _0955_ _2152_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__a221oi_2
X_5377_ _2863_ _0848_ _2980_ _0849_ _2083_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__a221oi_1
X_4328_ _3078_ _0843_ _1043_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__o21ai_1
X_4259_ _0335_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6275__137 clknet_1_0__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__2725_ clknet_0__2725_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2725_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3630_ _2902_ _2910_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3561_ _3109_ vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5300_ _1996_ _2000_ _2004_ _2007_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3492_ _3039_ _3040_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__nand2_1
X_5231_ _2800_ _0782_ _0841_ _0781_ _1938_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__a221oi_1
X_5162_ _2987_ _0872_ _0742_ _0873_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__a221oi_1
X_4113_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__clkbuf_8
X_5093_ _1801_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__nor2_1
X_4044_ _0419_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _0762_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5995_ _2481_ _2499_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1
+ vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__o21ai_1
X_4946_ _3143_ _3126_ _0336_ _3123_ _1656_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__a221oi_1
X_4877_ egd_top.BitStream_buffer.BS_buffer\[74\] _0930_ _0931_ egd_top.BitStream_buffer.BS_buffer\[77\]
+ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3828_ _0546_ _3084_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3759_ _2903_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__nand2_1
X_6478_ net220 _0311_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_5429_ _2125_ _2128_ _2132_ _2135_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4800_ _0551_ _0840_ _0412_ _0842_ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5780_ net10 _3066_ _2376_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4731_ _0933_ _0607_ _0934_ _2904_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__a22o_1
X_4662_ _0802_ _2802_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__nand2_1
X_6401_ net143 _0234_ net52 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[55\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3613_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6258__121 clknet_1_0__leaf__2726_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
X_4593_ _0892_ _2859_ _0893_ _0926_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__a221oi_1
X_3544_ _3092_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__clkbuf_4
X_3475_ _2946_ _2961_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5214_ _1921_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5145_ _0412_ _0840_ _3007_ _0842_ _1853_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__a221oi_1
X_5076_ _1075_ _0969_ _3129_ _0971_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__o22ai_1
X_4027_ _0377_ _0343_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nand2_1
X_5978_ _2551_ _2511_ _2512_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__nand3_1
X_4929_ _3115_ _0863_ _0864_ egd_top.BitStream_buffer.BS_buffer\[56\] _1639_ vssd1
+ vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__a221oi_2
X_6306__166 clknet_1_1__leaf__2729_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__inv_2
X_6196__64 clknet_1_0__leaf__2721_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__inv_2
Xclkbuf_0__2727_ _2727_ vssd1 vssd1 vccd1 vccd1 clknet_0__2727_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__clkbuf_8
X_3191_ egd_top.BitStream_buffer.pc_reg\[0\] _2760_ vssd1 vssd1 vccd1 vccd1 _2761_
+ sky130_fd_sc_hd__or2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5901_ _2472_ _2477_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5832_ net5 _0894_ _2420_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5763_ _2381_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4714_ _2974_ _3126_ _0333_ _3123_ _1426_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__a221oi_1
X_5694_ _2343_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_6327__17 clknet_1_1__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__inv_2
XFILLER_0_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4645_ _0526_ _0446_ _0619_ _0449_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__o22ai_1
X_4576_ _1280_ _1283_ _1286_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__and4_1
X_3527_ _2870_ _2937_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__nand2_1
X_3458_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__buf_4
X_3389_ _2884_ _2937_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__and2_1
X_5128_ _1826_ _1829_ _1832_ _1836_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__and4_2
X_5059_ _1185_ _3131_ _3108_ _3135_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6175__45 clknet_1_0__leaf__2719_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__inv_2
X_4430_ _1143_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__nand2_1
XANTENNA_2 _0444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6190__59 clknet_1_0__leaf__2720_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__inv_2
X_4361_ _0378_ _3126_ _0341_ _3123_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__a221oi_2
X_6100_ _2664_ _2668_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3312_ _2849_ _2854_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__o21ai_1
X_4292_ _0919_ _0953_ _0980_ _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__and4_1
X_3243_ net4 _2804_ _2798_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__mux2_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _2543_ _2457_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__nand2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ net29 vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__inv_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5815_ net36 egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5746_ _2798_ _2370_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5677_ egd_top.BitStream_buffer.buffer_index\[6\] _2795_ vssd1 vssd1 vccd1 vccd1
+ _2334_ sky130_fd_sc_hd__or2_4
XFILLER_0_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4628_ _0656_ _0961_ _0962_ _0371_ _1341_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4559_ _0833_ _2814_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__nand2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3930_ _0646_ _0647_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3861_ _0357_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0580_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3792_ _2997_ _2814_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand2_1
X_5600_ _2293_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
X_5531_ _3117_ _0366_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__nand2_1
X_5462_ _0791_ _2802_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4413_ _1115_ _1120_ _1124_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__and4_1
X_5393_ _0897_ _0926_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__nand2_1
X_4344_ _0874_ _0587_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__nand2_1
X_6014_ _2589_ _2552_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__nand2_1
X_4275_ _0424_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__clkbuf_4
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ net14 _0553_ _2353_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6252__116 clknet_1_0__leaf__2725_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _0777_ _0456_ _2789_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o21ai_1
X_4962_ _0904_ _0969_ _3108_ _0971_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__o22ai_1
X_4893_ _0797_ _2812_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__nand2_1
X_3913_ _2891_ _0629_ _0630_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3844_ _0560_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3775_ _0489_ _2945_ _0490_ _0491_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_54_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6311__2 clknet_1_1__leaf__2730_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__inv_2
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6494_ net68 egd_top.BitStream_buffer.pc\[2\] net36 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5514_ _0983_ _0882_ _2217_ _2218_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__o2111a_1
X_5445_ _0567_ _0956_ _1603_ _0958_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5376_ _0516_ _0850_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4327_ _0844_ _0443_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nand2_1
X_4258_ _0342_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__clkbuf_4
X_3209_ _2772_ _2777_ _2751_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4189_ _2935_ _3126_ _0378_ _3123_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2724_ clknet_0__2724_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2724_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3560_ _2893_ _2937_ vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__nand2_1
X_5230_ _0988_ _0783_ _0784_ _1116_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__a22o_1
X_3491_ egd_top.BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__buf_4
X_5161_ _1868_ _1869_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ _0824_ _2863_ _0825_ _2920_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__a221oi_1
X_5092_ _3067_ _0446_ _3031_ _0449_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__o22ai_1
X_4043_ _0417_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _0761_
+ sky130_fd_sc_hd__nand2_1
X_5994_ _2566_ _2569_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__nand2_1
X_4945_ _1066_ _3131_ _0543_ _3135_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _0937_ _2957_ _0656_ _0938_ _1587_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__a221oi_2
X_3827_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3758_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6235__100 clknet_1_0__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
X_3689_ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__clkbuf_4
X_6477_ net219 _0310_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[122\]
+ sky130_fd_sc_hd__dfrtp_2
X_5428_ _2133_ _2134_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__nor2_1
X_5359_ _3144_ _0811_ _2065_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4730_ egd_top.BitStream_buffer.BS_buffer\[73\] _0930_ _0931_ egd_top.BitStream_buffer.BS_buffer\[76\]
+ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ _1372_ _3065_ _0698_ _0796_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__o221a_1
X_6400_ net142 _0233_ net52 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[56\]
+ sky130_fd_sc_hd__dfrtp_4
X_3612_ _3156_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4592_ _1304_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__nand2_1
X_3543_ _2767_ _2865_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3474_ _3022_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _3023_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5213_ _0949_ _0656_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__nand2_1
X_5144_ _0516_ _0843_ _1852_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__o21ai_1
X_5075_ _2859_ _0961_ _0962_ _0709_ _1784_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__a221oi_1
X_4026_ _0741_ _0743_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5977_ net17 _2759_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__nor2_2
X_4928_ _1637_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2726_ _2726_ vssd1 vssd1 vccd1 vccd1 clknet_0__2726_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4859_ _0999_ _0587_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _2758_ _2759_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5900_ _2476_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5831_ _2422_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
X_5762_ net4 _2987_ _2377_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4713_ _0653_ _3131_ _0730_ _3135_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5693_ net15 egd_top.BitStream_buffer.BS_buffer\[55\] _2335_ vssd1 vssd1 vccd1 vccd1
+ _2343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4644_ _0439_ _0638_ _0441_ _0610_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4575_ _2907_ _0857_ _3127_ _0858_ _1288_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__a221oi_1
X_3526_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3457_ _2998_ _3000_ _3003_ _3005_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__and4_1
X_3388_ _2769_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__clkbuf_4
X_5127_ _2806_ _0800_ _0801_ _2828_ _1835_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5058_ _1724_ _1738_ _1750_ _1767_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__and4_1
X_4009_ _0337_ _0335_ _3133_ _0338_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 _0477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _1075_ _3131_ _0970_ _3135_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3311_ _2858_ _2859_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__nand2_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _0986_ _0995_ _1003_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__and4_1
X_3242_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__buf_4
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _2599_ _2509_ _2604_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__nand3_1
X_3173_ net28 vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__inv_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5814_ _2413_ _2401_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[3\] sky130_fd_sc_hd__xnor2_4
XFILLER_0_91_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5745_ _2795_ _2773_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5676_ _2333_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4627_ _0731_ _0963_ _0347_ _0964_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4558_ _0824_ _2913_ _0825_ _2980_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3509_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__clkbuf_8
X_4489_ _3087_ _0385_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__nand2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _0566_ _0570_ _0573_ _0578_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3791_ _0506_ _2982_ _0507_ _0508_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5530_ _2224_ _2228_ _2232_ _2235_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5461_ _2804_ _0782_ _0551_ _0781_ _2166_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4412_ _1125_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5392_ _0895_ _0469_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4343_ egd_top.BitStream_buffer.BS_buffer\[53\] _0863_ _0864_ _3112_ _1058_ vssd1
+ vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__a221oi_2
X_4274_ _0990_ _0477_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__nand2_1
X_6013_ _2588_ _2512_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__nand2_1
X_3225_ _2790_ _2782_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__nor2_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3989_ _3096_ _2907_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nand2_1
X_5728_ _2361_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5659_ net15 _0343_ _2317_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__mux2_1
X_6232__97 clknet_1_1__leaf__2724_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
XFILLER_0_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _0709_ _0961_ _0962_ _0553_ _1671_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__a221oi_1
X_4892_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3912_ _2866_ _2922_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3843_ _0561_ _3131_ _0349_ _3135_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3774_ _0492_ _2953_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__or2_1
X_6493_ net67 egd_top.BitStream_buffer.pc\[1\] net37 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5513_ _0889_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _2219_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5444_ _2139_ _2142_ _2146_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5375_ _2866_ _0341_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__nand2_1
X_4326_ _1031_ _1035_ _1037_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4257_ _0340_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__clkbuf_4
X_4188_ _0904_ _3131_ _0731_ _3135_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__o22ai_1
X_3208_ _2753_ _2776_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2777_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2723_ clknet_0__2723_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2723_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3490_ _2870_ _2915_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5160_ _0877_ _3112_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__nand2_1
X_4111_ _0407_ _0826_ _0757_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__o22ai_1
X_5091_ _0439_ _3034_ _0441_ _3048_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__a22o_1
X_4042_ _0758_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _2567_ _2568_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4944_ _1610_ _1624_ _1636_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__and4_1
XFILLER_0_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4875_ _1585_ _1586_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6211__78 clknet_1_1__leaf__2722_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
X_3826_ _0544_ _3080_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3757_ _2900_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _0476_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3688_ _2933_ _2915_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__nand2_1
X_6476_ net218 _0309_ net45 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[123\]
+ sky130_fd_sc_hd__dfrtp_2
X_5427_ _1533_ _3130_ _0717_ _3134_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__o22ai_1
X_5358_ _0812_ _3090_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__nand2_1
X_4309_ _0804_ _2822_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__nand2_1
X_5289_ _0990_ _3037_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6281__143 clknet_1_1__leaf__2727_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4660_ _0797_ _2808_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3611_ _2791_ _3157_ _0329_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4591_ _0897_ _0464_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__nand2_1
X_3542_ _3090_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3473_ _2927_ _2852_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__and2_1
X_6192_ clknet_1_0__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__buf_1
X_5212_ _0947_ _2957_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5143_ _0844_ _3053_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__nand2_1
X_5074_ _0730_ _0963_ _0543_ _0964_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ _0373_ egd_top.BitStream_buffer.BS_buffer\[88\] _0374_ _0742_ vssd1 vssd1
+ vccd1 vccd1 _0743_ sky130_fd_sc_hd__a22o_1
X_5976_ _2552_ _2513_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__nand2_1
X_4927_ _0867_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _1638_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2725_ _2725_ vssd1 vssd1 vccd1 vccd1 clknet_0__2725_ sky130_fd_sc_hd__clkbuf_16
X_4858_ _0428_ _0830_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__nand2_1
X_3809_ _3036_ _3053_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__nand2_1
X_4789_ _1499_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6459_ net201 _0292_ net38 vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6288__149 clknet_1_0__leaf__2728_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__inv_2
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5830_ net6 _0657_ _2420_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5761_ _2380_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4712_ _1379_ _1393_ _1406_ _1424_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__and4_1
X_5692_ _2342_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4643_ _0709_ _0996_ _0463_ _0997_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__a221oi_1
X_4574_ _1287_ _2912_ _0641_ _2917_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3525_ _2925_ _2979_ _3029_ _3073_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__and4_1
X_6244_ clknet_1_1__leaf__2717_ vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__buf_1
X_3456_ _3004_ _2804_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__nand2_1
X_3387_ _2934_ _2935_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5126_ _1833_ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__nand2_1
X_5057_ _1754_ _1758_ _1762_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4008_ _0724_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5959_ _2530_ _2535_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_4 _0477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3310_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__buf_4
X_6332__22 clknet_1_0__leaf__2731_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__inv_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _1004_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__nor2_1
X_3241_ _2803_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__clkbuf_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ net30 vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__inv_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5813_ _2402_ _2403_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ _2369_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5675_ net1 _2931_ _2316_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4626_ _2810_ _0954_ _2808_ _0955_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_32_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4557_ _0984_ _0826_ _0601_ _0827_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__o22ai_1
X_3508_ _2833_ _2985_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__and2_1
X_4488_ _0489_ _3084_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__or2_1
X_3439_ _2986_ _2987_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__nand2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _1807_ _1811_ _1815_ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__and4_1
X_6089_ _2653_ _2554_ _2658_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__nand3_1
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 la_data_out_18_16[2] sky130_fd_sc_hd__buf_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _2992_ _3010_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__nand2_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5460_ _0841_ _0783_ _0784_ _3101_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4411_ _1126_ _0446_ _3151_ _0449_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5391_ _3048_ _0872_ _0871_ _0873_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4342_ _1056_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__nand2_1
X_4273_ _0419_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__buf_4
X_6012_ _2575_ _2587_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__nand2_1
X_3224_ _2789_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__clkbuf_4
.ends

