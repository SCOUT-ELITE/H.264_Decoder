// This is the unpowered netlist.
module egd_top_wrapper (wb_clk_i,
    wb_rst_i,
    la_data_in_47_32,
    la_data_in_49_48,
    la_data_out_15_8,
    la_data_out_18_16,
    la_data_out_22_19);
 input wb_clk_i;
 input wb_rst_i;
 input [15:0] la_data_in_47_32;
 input [1:0] la_data_in_49_48;
 output [7:0] la_data_out_15_8;
 output [2:0] la_data_out_18_16;
 output [3:0] la_data_out_22_19;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire \egd_top.BitStream_buffer.BS_buffer[0] ;
 wire \egd_top.BitStream_buffer.BS_buffer[100] ;
 wire \egd_top.BitStream_buffer.BS_buffer[101] ;
 wire \egd_top.BitStream_buffer.BS_buffer[102] ;
 wire \egd_top.BitStream_buffer.BS_buffer[103] ;
 wire \egd_top.BitStream_buffer.BS_buffer[104] ;
 wire \egd_top.BitStream_buffer.BS_buffer[105] ;
 wire \egd_top.BitStream_buffer.BS_buffer[106] ;
 wire \egd_top.BitStream_buffer.BS_buffer[107] ;
 wire \egd_top.BitStream_buffer.BS_buffer[108] ;
 wire \egd_top.BitStream_buffer.BS_buffer[109] ;
 wire \egd_top.BitStream_buffer.BS_buffer[10] ;
 wire \egd_top.BitStream_buffer.BS_buffer[110] ;
 wire \egd_top.BitStream_buffer.BS_buffer[111] ;
 wire \egd_top.BitStream_buffer.BS_buffer[112] ;
 wire \egd_top.BitStream_buffer.BS_buffer[113] ;
 wire \egd_top.BitStream_buffer.BS_buffer[114] ;
 wire \egd_top.BitStream_buffer.BS_buffer[115] ;
 wire \egd_top.BitStream_buffer.BS_buffer[116] ;
 wire \egd_top.BitStream_buffer.BS_buffer[117] ;
 wire \egd_top.BitStream_buffer.BS_buffer[118] ;
 wire \egd_top.BitStream_buffer.BS_buffer[119] ;
 wire \egd_top.BitStream_buffer.BS_buffer[11] ;
 wire \egd_top.BitStream_buffer.BS_buffer[120] ;
 wire \egd_top.BitStream_buffer.BS_buffer[121] ;
 wire \egd_top.BitStream_buffer.BS_buffer[122] ;
 wire \egd_top.BitStream_buffer.BS_buffer[123] ;
 wire \egd_top.BitStream_buffer.BS_buffer[124] ;
 wire \egd_top.BitStream_buffer.BS_buffer[125] ;
 wire \egd_top.BitStream_buffer.BS_buffer[126] ;
 wire \egd_top.BitStream_buffer.BS_buffer[127] ;
 wire \egd_top.BitStream_buffer.BS_buffer[12] ;
 wire \egd_top.BitStream_buffer.BS_buffer[13] ;
 wire \egd_top.BitStream_buffer.BS_buffer[14] ;
 wire \egd_top.BitStream_buffer.BS_buffer[15] ;
 wire \egd_top.BitStream_buffer.BS_buffer[16] ;
 wire \egd_top.BitStream_buffer.BS_buffer[17] ;
 wire \egd_top.BitStream_buffer.BS_buffer[18] ;
 wire \egd_top.BitStream_buffer.BS_buffer[19] ;
 wire \egd_top.BitStream_buffer.BS_buffer[1] ;
 wire \egd_top.BitStream_buffer.BS_buffer[20] ;
 wire \egd_top.BitStream_buffer.BS_buffer[21] ;
 wire \egd_top.BitStream_buffer.BS_buffer[22] ;
 wire \egd_top.BitStream_buffer.BS_buffer[23] ;
 wire \egd_top.BitStream_buffer.BS_buffer[24] ;
 wire \egd_top.BitStream_buffer.BS_buffer[25] ;
 wire \egd_top.BitStream_buffer.BS_buffer[26] ;
 wire \egd_top.BitStream_buffer.BS_buffer[27] ;
 wire \egd_top.BitStream_buffer.BS_buffer[28] ;
 wire \egd_top.BitStream_buffer.BS_buffer[29] ;
 wire \egd_top.BitStream_buffer.BS_buffer[2] ;
 wire \egd_top.BitStream_buffer.BS_buffer[30] ;
 wire \egd_top.BitStream_buffer.BS_buffer[31] ;
 wire \egd_top.BitStream_buffer.BS_buffer[32] ;
 wire \egd_top.BitStream_buffer.BS_buffer[33] ;
 wire \egd_top.BitStream_buffer.BS_buffer[34] ;
 wire \egd_top.BitStream_buffer.BS_buffer[35] ;
 wire \egd_top.BitStream_buffer.BS_buffer[36] ;
 wire \egd_top.BitStream_buffer.BS_buffer[37] ;
 wire \egd_top.BitStream_buffer.BS_buffer[38] ;
 wire \egd_top.BitStream_buffer.BS_buffer[39] ;
 wire \egd_top.BitStream_buffer.BS_buffer[3] ;
 wire \egd_top.BitStream_buffer.BS_buffer[40] ;
 wire \egd_top.BitStream_buffer.BS_buffer[41] ;
 wire \egd_top.BitStream_buffer.BS_buffer[42] ;
 wire \egd_top.BitStream_buffer.BS_buffer[43] ;
 wire \egd_top.BitStream_buffer.BS_buffer[44] ;
 wire \egd_top.BitStream_buffer.BS_buffer[45] ;
 wire \egd_top.BitStream_buffer.BS_buffer[46] ;
 wire \egd_top.BitStream_buffer.BS_buffer[47] ;
 wire \egd_top.BitStream_buffer.BS_buffer[48] ;
 wire \egd_top.BitStream_buffer.BS_buffer[49] ;
 wire \egd_top.BitStream_buffer.BS_buffer[4] ;
 wire \egd_top.BitStream_buffer.BS_buffer[50] ;
 wire \egd_top.BitStream_buffer.BS_buffer[51] ;
 wire \egd_top.BitStream_buffer.BS_buffer[52] ;
 wire \egd_top.BitStream_buffer.BS_buffer[53] ;
 wire \egd_top.BitStream_buffer.BS_buffer[54] ;
 wire \egd_top.BitStream_buffer.BS_buffer[55] ;
 wire \egd_top.BitStream_buffer.BS_buffer[56] ;
 wire \egd_top.BitStream_buffer.BS_buffer[57] ;
 wire \egd_top.BitStream_buffer.BS_buffer[58] ;
 wire \egd_top.BitStream_buffer.BS_buffer[59] ;
 wire \egd_top.BitStream_buffer.BS_buffer[5] ;
 wire \egd_top.BitStream_buffer.BS_buffer[60] ;
 wire \egd_top.BitStream_buffer.BS_buffer[61] ;
 wire \egd_top.BitStream_buffer.BS_buffer[62] ;
 wire \egd_top.BitStream_buffer.BS_buffer[63] ;
 wire \egd_top.BitStream_buffer.BS_buffer[64] ;
 wire \egd_top.BitStream_buffer.BS_buffer[65] ;
 wire \egd_top.BitStream_buffer.BS_buffer[66] ;
 wire \egd_top.BitStream_buffer.BS_buffer[67] ;
 wire \egd_top.BitStream_buffer.BS_buffer[68] ;
 wire \egd_top.BitStream_buffer.BS_buffer[69] ;
 wire \egd_top.BitStream_buffer.BS_buffer[6] ;
 wire \egd_top.BitStream_buffer.BS_buffer[70] ;
 wire \egd_top.BitStream_buffer.BS_buffer[71] ;
 wire \egd_top.BitStream_buffer.BS_buffer[72] ;
 wire \egd_top.BitStream_buffer.BS_buffer[73] ;
 wire \egd_top.BitStream_buffer.BS_buffer[74] ;
 wire \egd_top.BitStream_buffer.BS_buffer[75] ;
 wire \egd_top.BitStream_buffer.BS_buffer[76] ;
 wire \egd_top.BitStream_buffer.BS_buffer[77] ;
 wire \egd_top.BitStream_buffer.BS_buffer[78] ;
 wire \egd_top.BitStream_buffer.BS_buffer[79] ;
 wire \egd_top.BitStream_buffer.BS_buffer[7] ;
 wire \egd_top.BitStream_buffer.BS_buffer[80] ;
 wire \egd_top.BitStream_buffer.BS_buffer[81] ;
 wire \egd_top.BitStream_buffer.BS_buffer[82] ;
 wire \egd_top.BitStream_buffer.BS_buffer[83] ;
 wire \egd_top.BitStream_buffer.BS_buffer[84] ;
 wire \egd_top.BitStream_buffer.BS_buffer[85] ;
 wire \egd_top.BitStream_buffer.BS_buffer[86] ;
 wire \egd_top.BitStream_buffer.BS_buffer[87] ;
 wire \egd_top.BitStream_buffer.BS_buffer[88] ;
 wire \egd_top.BitStream_buffer.BS_buffer[89] ;
 wire \egd_top.BitStream_buffer.BS_buffer[8] ;
 wire \egd_top.BitStream_buffer.BS_buffer[90] ;
 wire \egd_top.BitStream_buffer.BS_buffer[91] ;
 wire \egd_top.BitStream_buffer.BS_buffer[92] ;
 wire \egd_top.BitStream_buffer.BS_buffer[93] ;
 wire \egd_top.BitStream_buffer.BS_buffer[94] ;
 wire \egd_top.BitStream_buffer.BS_buffer[95] ;
 wire \egd_top.BitStream_buffer.BS_buffer[96] ;
 wire \egd_top.BitStream_buffer.BS_buffer[97] ;
 wire \egd_top.BitStream_buffer.BS_buffer[98] ;
 wire \egd_top.BitStream_buffer.BS_buffer[99] ;
 wire \egd_top.BitStream_buffer.BS_buffer[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[10] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[11] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[12] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[13] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[14] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[15] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[1] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[2] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[3] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[4] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[5] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[6] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[7] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[8] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_valid_n ;
 wire \egd_top.BitStream_buffer.buffer_index[4] ;
 wire \egd_top.BitStream_buffer.buffer_index[5] ;
 wire \egd_top.BitStream_buffer.buffer_index[6] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[1] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[2] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[3] ;
 wire \egd_top.BitStream_buffer.pc[0] ;
 wire \egd_top.BitStream_buffer.pc[1] ;
 wire \egd_top.BitStream_buffer.pc[2] ;
 wire \egd_top.BitStream_buffer.pc[3] ;
 wire \egd_top.BitStream_buffer.pc[4] ;
 wire \egd_top.BitStream_buffer.pc[5] ;
 wire \egd_top.BitStream_buffer.pc[6] ;
 wire \egd_top.BitStream_buffer.pc_previous[0] ;
 wire \egd_top.BitStream_buffer.pc_previous[1] ;
 wire \egd_top.BitStream_buffer.pc_previous[2] ;
 wire \egd_top.BitStream_buffer.pc_previous[3] ;
 wire \egd_top.BitStream_buffer.pc_previous[4] ;
 wire \egd_top.BitStream_buffer.pc_previous[5] ;
 wire \egd_top.BitStream_buffer.pc_previous[6] ;
 wire \egd_top.BitStream_buffer.pc_reg[0] ;
 wire \egd_top.BitStream_buffer.pc_reg[1] ;
 wire \egd_top.BitStream_buffer.pc_reg[2] ;
 wire \egd_top.BitStream_buffer.pc_reg[3] ;
 wire \egd_top.BitStream_buffer.pc_reg[4] ;
 wire \egd_top.BitStream_buffer.pc_reg[5] ;
 wire \egd_top.BitStream_buffer.pc_reg[6] ;
 wire \egd_top.exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_1855_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_1972_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_2269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_2269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_2821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_2859_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_3104_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_2900_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0889_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1514_));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_91 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3152_ (.A(net33),
    .Y(_2718_));
 sky130_fd_sc_hd__nand2_1 _3153_ (.A(net32),
    .B(net31),
    .Y(_2719_));
 sky130_fd_sc_hd__inv_2 _3154_ (.A(net34),
    .Y(_2720_));
 sky130_fd_sc_hd__o21ai_1 _3155_ (.A1(_2718_),
    .A2(_2719_),
    .B1(_2720_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor2_1 _3156_ (.A(net33),
    .B(net32),
    .Y(_2721_));
 sky130_fd_sc_hd__nor2_1 _3157_ (.A(_2720_),
    .B(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__inv_2 _3158_ (.A(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__a21o_1 _3159_ (.A1(_2718_),
    .A2(_2719_),
    .B1(_0321_),
    .X(_2724_));
 sky130_fd_sc_hd__o21ai_1 _3160_ (.A1(_2718_),
    .A2(_2723_),
    .B1(_2724_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _3161_ (.A(net31),
    .Y(_2725_));
 sky130_fd_sc_hd__nor2_1 _3162_ (.A(_2725_),
    .B(_2722_),
    .Y(_2726_));
 sky130_fd_sc_hd__o22a_1 _3163_ (.A1(_2719_),
    .A2(_2722_),
    .B1(net32),
    .B2(_2726_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_1 _3164_ (.A(net31),
    .B(_2723_),
    .Y(_2727_));
 sky130_fd_sc_hd__nor2_1 _3165_ (.A(_2726_),
    .B(_2727_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _3166_ (.A(net30),
    .Y(_2728_));
 sky130_fd_sc_hd__inv_2 _3167_ (.A(net28),
    .Y(_2729_));
 sky130_fd_sc_hd__inv_2 _3168_ (.A(net29),
    .Y(_2730_));
 sky130_fd_sc_hd__nand2_1 _3169_ (.A(_2728_),
    .B(_2730_),
    .Y(_2731_));
 sky130_fd_sc_hd__nand2_1 _3170_ (.A(_2729_),
    .B(net29),
    .Y(_2732_));
 sky130_fd_sc_hd__o211a_1 _3171_ (.A1(_2728_),
    .A2(_2729_),
    .B1(_2731_),
    .C1(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__nand2_1 _3172_ (.A(_2730_),
    .B(net28),
    .Y(_2734_));
 sky130_fd_sc_hd__nand2_1 _3173_ (.A(net30),
    .B(net29),
    .Y(_2735_));
 sky130_fd_sc_hd__nor2_1 _3174_ (.A(net28),
    .B(_2731_),
    .Y(_2736_));
 sky130_fd_sc_hd__inv_2 _3175_ (.A(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__o211ai_2 _3176_ (.A1(_2728_),
    .A2(_2734_),
    .B1(_2735_),
    .C1(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__nand2_1 _3177_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_2739_));
 sky130_fd_sc_hd__nand2_1 _3178_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.pc_previous[2] ),
    .Y(_2740_));
 sky130_fd_sc_hd__nand2_1 _3179_ (.A(\egd_top.BitStream_buffer.pc_previous[5] ),
    .B(\egd_top.BitStream_buffer.pc_previous[4] ),
    .Y(_2741_));
 sky130_fd_sc_hd__or3_1 _3180_ (.A(_2739_),
    .B(_2740_),
    .C(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__inv_2 _3181_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .Y(_2743_));
 sky130_fd_sc_hd__nand2_4 _3182_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .B(net39),
    .Y(_2744_));
 sky130_fd_sc_hd__inv_2 _3183_ (.A(net17),
    .Y(_2745_));
 sky130_fd_sc_hd__inv_2 _3184_ (.A(net18),
    .Y(_2746_));
 sky130_fd_sc_hd__nand2_1 _3185_ (.A(_2745_),
    .B(_2746_),
    .Y(_2747_));
 sky130_fd_sc_hd__or2_1 _3186_ (.A(\egd_top.BitStream_buffer.pc_reg[0] ),
    .B(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__buf_6 _3187_ (.A(_2747_),
    .X(_2749_));
 sky130_fd_sc_hd__nand2_4 _3188_ (.A(_2749_),
    .B(\egd_top.BitStream_buffer.pc_reg[0] ),
    .Y(_2750_));
 sky130_fd_sc_hd__nand2_4 _3189_ (.A(_2748_),
    .B(_2750_),
    .Y(_2751_));
 sky130_fd_sc_hd__clkinv_4 _3190_ (.A(_2751_),
    .Y(\egd_top.BitStream_buffer.pc[0] ));
 sky130_fd_sc_hd__nand2_4 _3191_ (.A(\egd_top.BitStream_buffer.pc[0] ),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2752_));
 sky130_fd_sc_hd__nor2_4 _3192_ (.A(_2744_),
    .B(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__inv_2 _3193_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2754_));
 sky130_fd_sc_hd__and3_2 _3194_ (.A(_2754_),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_2755_));
 sky130_fd_sc_hd__and2_1 _3195_ (.A(_2753_),
    .B(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__buf_2 _3196_ (.A(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__a211o_1 _3197_ (.A1(_2742_),
    .A2(_2743_),
    .B1(\egd_top.BitStream_buffer.pc[6] ),
    .C1(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__inv_2 _3198_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .Y(_2759_));
 sky130_fd_sc_hd__inv_2 _3199_ (.A(\egd_top.BitStream_buffer.buffer_index[5] ),
    .Y(_2760_));
 sky130_fd_sc_hd__inv_2 _3200_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_2761_));
 sky130_fd_sc_hd__and3_1 _3201_ (.A(_2759_),
    .B(_2760_),
    .C(_2761_),
    .X(_2762_));
 sky130_fd_sc_hd__o21ai_1 _3202_ (.A1(_2743_),
    .A2(_2762_),
    .B1(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2763_));
 sky130_fd_sc_hd__a21o_1 _3203_ (.A1(_2758_),
    .A2(_2763_),
    .B1(_2737_),
    .X(_2764_));
 sky130_fd_sc_hd__and3_1 _3204_ (.A(_2760_),
    .B(_2761_),
    .C(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(_2765_));
 sky130_fd_sc_hd__or4b_1 _3205_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_2737_),
    .C(_2757_),
    .D_N(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__o2111ai_1 _3206_ (.A1(_2728_),
    .A2(_2734_),
    .B1(_2738_),
    .C1(_2764_),
    .D1(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__and4_1 _3207_ (.A(_2718_),
    .B(_2725_),
    .C(net34),
    .D(net32),
    .X(_2768_));
 sky130_fd_sc_hd__nand2_1 _3208_ (.A(_2767_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(_2733_),
    .A1(net30),
    .S(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_2770_),
    .X(_0317_));
 sky130_fd_sc_hd__a21oi_1 _3211_ (.A1(_2734_),
    .A2(_2732_),
    .B1(net30),
    .Y(_2771_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(_2771_),
    .A1(net29),
    .S(_2769_),
    .X(_2772_));
 sky130_fd_sc_hd__clkbuf_1 _3213_ (.A(_2772_),
    .X(_0316_));
 sky130_fd_sc_hd__o211ai_1 _3214_ (.A1(net28),
    .A2(_2738_),
    .B1(_2764_),
    .C1(_2766_),
    .Y(_2773_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(_2773_),
    .A1(net28),
    .S(_2769_),
    .X(_2774_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_2774_),
    .X(_0315_));
 sky130_fd_sc_hd__inv_2 _3217_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .Y(_2775_));
 sky130_fd_sc_hd__clkbuf_4 _3218_ (.A(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__nor2_1 _3219_ (.A(_2776_),
    .B(_2768_),
    .Y(_0314_));
 sky130_fd_sc_hd__buf_4 _3220_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .X(_2777_));
 sky130_fd_sc_hd__nand2_1 _3221_ (.A(_2721_),
    .B(_2720_),
    .Y(_2778_));
 sky130_fd_sc_hd__a22o_2 _3222_ (.A1(_2731_),
    .A2(_2735_),
    .B1(_2723_),
    .B2(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__nand2_1 _3223_ (.A(_2779_),
    .B(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_2780_));
 sky130_fd_sc_hd__or2_1 _3224_ (.A(_2760_),
    .B(_2780_),
    .X(_2781_));
 sky130_fd_sc_hd__or2_1 _3225_ (.A(_2759_),
    .B(_2781_),
    .X(_2782_));
 sky130_fd_sc_hd__buf_2 _3226_ (.A(_2782_),
    .X(_2783_));
 sky130_fd_sc_hd__buf_4 _3227_ (.A(_2783_),
    .X(_2784_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(net7),
    .A1(_2777_),
    .S(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__clkbuf_1 _3229_ (.A(_2785_),
    .X(_0313_));
 sky130_fd_sc_hd__buf_4 _3230_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_2786_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(net6),
    .A1(_2786_),
    .S(_2784_),
    .X(_2787_));
 sky130_fd_sc_hd__clkbuf_1 _3232_ (.A(_2787_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_4 _3233_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .X(_2788_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(net5),
    .A1(_2788_),
    .S(_2784_),
    .X(_2789_));
 sky130_fd_sc_hd__clkbuf_1 _3235_ (.A(_2789_),
    .X(_0311_));
 sky130_fd_sc_hd__buf_4 _3236_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .X(_2790_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(net4),
    .A1(_2790_),
    .S(_2784_),
    .X(_2791_));
 sky130_fd_sc_hd__clkbuf_1 _3238_ (.A(_2791_),
    .X(_0310_));
 sky130_fd_sc_hd__buf_4 _3239_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .X(_2792_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(net3),
    .A1(_2792_),
    .S(_2784_),
    .X(_2793_));
 sky130_fd_sc_hd__clkbuf_1 _3241_ (.A(_2793_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_4 _3242_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .X(_2794_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(net2),
    .A1(_2794_),
    .S(_2784_),
    .X(_2795_));
 sky130_fd_sc_hd__clkbuf_1 _3244_ (.A(_2795_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_4 _3245_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .X(_2796_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(net16),
    .A1(_2796_),
    .S(_2784_),
    .X(_2797_));
 sky130_fd_sc_hd__clkbuf_1 _3247_ (.A(_2797_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_4 _3248_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_2798_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(net15),
    .A1(_2798_),
    .S(_2784_),
    .X(_2799_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_2799_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_4 _3251_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_2800_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(net14),
    .A1(_2800_),
    .S(_2784_),
    .X(_2801_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_2801_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_4 _3254_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_2802_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(net13),
    .A1(_2802_),
    .S(_2784_),
    .X(_2803_));
 sky130_fd_sc_hd__clkbuf_1 _3256_ (.A(_2803_),
    .X(_0304_));
 sky130_fd_sc_hd__buf_4 _3257_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_2804_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(net12),
    .A1(_2804_),
    .S(_2784_),
    .X(_2805_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_2805_),
    .X(_0303_));
 sky130_fd_sc_hd__buf_4 _3260_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .X(_2806_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(net11),
    .A1(_2806_),
    .S(_2783_),
    .X(_2807_));
 sky130_fd_sc_hd__clkbuf_1 _3262_ (.A(_2807_),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_8 _3263_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_2808_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(net10),
    .A1(_2808_),
    .S(_2783_),
    .X(_2809_));
 sky130_fd_sc_hd__clkbuf_1 _3265_ (.A(_2809_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_8 _3266_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_2810_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(net9),
    .A1(_2810_),
    .S(_2783_),
    .X(_2811_));
 sky130_fd_sc_hd__clkbuf_1 _3268_ (.A(_2811_),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_8 _3269_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_2812_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(net8),
    .A1(_2812_),
    .S(_2783_),
    .X(_2813_));
 sky130_fd_sc_hd__clkbuf_1 _3271_ (.A(_2813_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_4 _3272_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_2814_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(net1),
    .A1(_2814_),
    .S(_2783_),
    .X(_2815_));
 sky130_fd_sc_hd__clkbuf_1 _3274_ (.A(_2815_),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_4 _3275_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .X(_2816_));
 sky130_fd_sc_hd__clkbuf_8 _3276_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_2817_));
 sky130_fd_sc_hd__inv_4 _3277_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_2818_));
 sky130_fd_sc_hd__inv_2 _3278_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2819_));
 sky130_fd_sc_hd__nand2_4 _3279_ (.A(_2751_),
    .B(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__nor3_4 _3280_ (.A(_2818_),
    .B(net39),
    .C(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__inv_2 _3281_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_2822_));
 sky130_fd_sc_hd__or3_1 _3282_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .B(_2754_),
    .C(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__inv_2 _3283_ (.A(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__and2_1 _3284_ (.A(_2821_),
    .B(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__clkbuf_2 _3285_ (.A(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__buf_4 _3286_ (.A(_2826_),
    .X(_2827_));
 sky130_fd_sc_hd__clkbuf_8 _3287_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_2828_));
 sky130_fd_sc_hd__nor3_2 _3288_ (.A(_2818_),
    .B(net39),
    .C(_2752_),
    .Y(_2829_));
 sky130_fd_sc_hd__and2_1 _3289_ (.A(net37),
    .B(_2824_),
    .X(_2830_));
 sky130_fd_sc_hd__clkbuf_2 _3290_ (.A(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__buf_4 _3291_ (.A(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__nand2_8 _3292_ (.A(\egd_top.BitStream_buffer.pc[0] ),
    .B(_2819_),
    .Y(_2833_));
 sky130_fd_sc_hd__nor3_4 _3293_ (.A(_2818_),
    .B(net39),
    .C(_2833_),
    .Y(_2834_));
 sky130_fd_sc_hd__and3_2 _3294_ (.A(_2754_),
    .B(_2822_),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_2835_));
 sky130_fd_sc_hd__clkbuf_4 _3295_ (.A(_2835_),
    .X(_2836_));
 sky130_fd_sc_hd__and2_1 _3296_ (.A(net36),
    .B(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__buf_4 _3297_ (.A(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__buf_4 _3298_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .X(_2839_));
 sky130_fd_sc_hd__nand2_1 _3299_ (.A(_2838_),
    .B(_2839_),
    .Y(_2840_));
 sky130_fd_sc_hd__nand2_8 _3300_ (.A(_2818_),
    .B(net39),
    .Y(_2841_));
 sky130_fd_sc_hd__nor2_8 _3301_ (.A(_2841_),
    .B(_2820_),
    .Y(_2842_));
 sky130_fd_sc_hd__clkbuf_4 _3302_ (.A(_2824_),
    .X(_2843_));
 sky130_fd_sc_hd__and2_1 _3303_ (.A(_2842_),
    .B(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__clkbuf_4 _3304_ (.A(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__clkbuf_8 _3305_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .X(_2846_));
 sky130_fd_sc_hd__nand2_1 _3306_ (.A(_2845_),
    .B(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__nand2_1 _3307_ (.A(_2840_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__a221oi_2 _3308_ (.A1(_2817_),
    .A2(_2827_),
    .B1(_2828_),
    .B2(_2832_),
    .C1(_2848_),
    .Y(_2849_));
 sky130_fd_sc_hd__nor2_4 _3309_ (.A(_2744_),
    .B(_2820_),
    .Y(_2850_));
 sky130_fd_sc_hd__and3_1 _3310_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_2851_));
 sky130_fd_sc_hd__buf_2 _3311_ (.A(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__and2_1 _3312_ (.A(_2850_),
    .B(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__clkbuf_4 _3313_ (.A(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__nor2_4 _3314_ (.A(_2841_),
    .B(_2752_),
    .Y(_2855_));
 sky130_fd_sc_hd__and2_1 _3315_ (.A(_2855_),
    .B(_2852_),
    .X(_2856_));
 sky130_fd_sc_hd__clkbuf_4 _3316_ (.A(_2856_),
    .X(_2857_));
 sky130_fd_sc_hd__a22o_1 _3317_ (.A1(_2854_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .B1(_2857_),
    .B2(_2806_),
    .X(_2858_));
 sky130_fd_sc_hd__nor2_4 _3318_ (.A(_2744_),
    .B(_2833_),
    .Y(_2859_));
 sky130_fd_sc_hd__clkbuf_4 _3319_ (.A(_2852_),
    .X(_2860_));
 sky130_fd_sc_hd__nand2_1 _3320_ (.A(_2859_),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__inv_2 _3321_ (.A(_2861_),
    .Y(_2862_));
 sky130_fd_sc_hd__nand2_1 _3322_ (.A(net36),
    .B(_2843_),
    .Y(_2863_));
 sky130_fd_sc_hd__inv_2 _3323_ (.A(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__clkbuf_8 _3324_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_2865_));
 sky130_fd_sc_hd__a22o_1 _3325_ (.A1(_2810_),
    .A2(_2862_),
    .B1(_2864_),
    .B2(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__nor2_1 _3326_ (.A(_2858_),
    .B(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__inv_2 _3327_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_2868_));
 sky130_fd_sc_hd__nand2_1 _3328_ (.A(_2850_),
    .B(_2843_),
    .Y(_2869_));
 sky130_fd_sc_hd__clkbuf_4 _3329_ (.A(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__inv_2 _3330_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_2871_));
 sky130_fd_sc_hd__inv_2 _3331_ (.A(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2872_));
 sky130_fd_sc_hd__nand2_4 _3332_ (.A(_2818_),
    .B(_2872_),
    .Y(_2873_));
 sky130_fd_sc_hd__nor2_8 _3333_ (.A(_2873_),
    .B(_2833_),
    .Y(_2874_));
 sky130_fd_sc_hd__nand2_4 _3334_ (.A(_2874_),
    .B(_2860_),
    .Y(_2875_));
 sky130_fd_sc_hd__nand2_4 _3335_ (.A(_2751_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2876_));
 sky130_fd_sc_hd__nor2_4 _3336_ (.A(_2744_),
    .B(_2876_),
    .Y(_2877_));
 sky130_fd_sc_hd__and2_1 _3337_ (.A(_2877_),
    .B(_2843_),
    .X(_2878_));
 sky130_fd_sc_hd__clkbuf_4 _3338_ (.A(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__buf_4 _3339_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .X(_2880_));
 sky130_fd_sc_hd__nand2_1 _3340_ (.A(_2879_),
    .B(_2880_),
    .Y(_2881_));
 sky130_fd_sc_hd__o221a_1 _3341_ (.A1(_2868_),
    .A2(_2870_),
    .B1(_2871_),
    .B2(_2875_),
    .C1(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__nor2_8 _3342_ (.A(_2841_),
    .B(_2833_),
    .Y(_2883_));
 sky130_fd_sc_hd__and2_1 _3343_ (.A(_2883_),
    .B(_2843_),
    .X(_2884_));
 sky130_fd_sc_hd__clkbuf_4 _3344_ (.A(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__clkbuf_8 _3345_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .X(_2886_));
 sky130_fd_sc_hd__and2_1 _3346_ (.A(_2821_),
    .B(_2860_),
    .X(_2887_));
 sky130_fd_sc_hd__clkbuf_4 _3347_ (.A(_2887_),
    .X(_2888_));
 sky130_fd_sc_hd__and2_1 _3348_ (.A(_2855_),
    .B(_2843_),
    .X(_2889_));
 sky130_fd_sc_hd__clkbuf_4 _3349_ (.A(_2889_),
    .X(_2890_));
 sky130_fd_sc_hd__clkbuf_8 _3350_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .X(_2891_));
 sky130_fd_sc_hd__nand2_1 _3351_ (.A(_2890_),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__and2_1 _3352_ (.A(_2842_),
    .B(_2860_),
    .X(_2893_));
 sky130_fd_sc_hd__clkbuf_4 _3353_ (.A(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__nand2_1 _3354_ (.A(_2894_),
    .B(_2800_),
    .Y(_2895_));
 sky130_fd_sc_hd__nand2_1 _3355_ (.A(_2892_),
    .B(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__a221oi_1 _3356_ (.A1(_2885_),
    .A2(_2886_),
    .B1(_2888_),
    .B2(_2792_),
    .C1(_2896_),
    .Y(_2897_));
 sky130_fd_sc_hd__and4_1 _3357_ (.A(_2849_),
    .B(_2867_),
    .C(_2882_),
    .D(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__buf_4 _3358_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .X(_2899_));
 sky130_fd_sc_hd__nor3_2 _3359_ (.A(_2818_),
    .B(net39),
    .C(_2876_),
    .Y(_2900_));
 sky130_fd_sc_hd__and2_1 _3360_ (.A(net35),
    .B(_2836_),
    .X(_2901_));
 sky130_fd_sc_hd__buf_1 _3361_ (.A(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__clkbuf_4 _3362_ (.A(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__clkbuf_8 _3363_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .X(_2904_));
 sky130_fd_sc_hd__and2_1 _3364_ (.A(net37),
    .B(_2836_),
    .X(_2905_));
 sky130_fd_sc_hd__buf_1 _3365_ (.A(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__buf_4 _3366_ (.A(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__buf_4 _3367_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .X(_2908_));
 sky130_fd_sc_hd__inv_2 _3368_ (.A(_2908_),
    .Y(_2909_));
 sky130_fd_sc_hd__nand2_1 _3369_ (.A(_2874_),
    .B(_2836_),
    .Y(_2910_));
 sky130_fd_sc_hd__clkbuf_4 _3370_ (.A(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__buf_6 _3371_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .X(_2912_));
 sky130_fd_sc_hd__clkinv_4 _3372_ (.A(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__nor2_4 _3373_ (.A(_2873_),
    .B(_2752_),
    .Y(_2914_));
 sky130_fd_sc_hd__nand2_1 _3374_ (.A(_2914_),
    .B(_2836_),
    .Y(_2915_));
 sky130_fd_sc_hd__clkbuf_4 _3375_ (.A(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__o22ai_1 _3376_ (.A1(_2909_),
    .A2(_2911_),
    .B1(_2913_),
    .B2(_2916_),
    .Y(_2917_));
 sky130_fd_sc_hd__a221oi_1 _3377_ (.A1(_2899_),
    .A2(_2903_),
    .B1(_2904_),
    .B2(_2907_),
    .C1(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__and2_1 _3378_ (.A(net35),
    .B(_2843_),
    .X(_2919_));
 sky130_fd_sc_hd__clkbuf_4 _3379_ (.A(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__clkbuf_8 _3380_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .X(_2921_));
 sky130_fd_sc_hd__and2_1 _3381_ (.A(net37),
    .B(_2860_),
    .X(_2922_));
 sky130_fd_sc_hd__clkbuf_4 _3382_ (.A(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__and2_1 _3383_ (.A(net35),
    .B(_2860_),
    .X(_2924_));
 sky130_fd_sc_hd__clkbuf_4 _3384_ (.A(_2924_),
    .X(_2925_));
 sky130_fd_sc_hd__nand2_1 _3385_ (.A(_2925_),
    .B(_2796_),
    .Y(_2926_));
 sky130_fd_sc_hd__and2_1 _3386_ (.A(_2914_),
    .B(_2860_),
    .X(_2927_));
 sky130_fd_sc_hd__clkbuf_4 _3387_ (.A(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__nand2_1 _3388_ (.A(_2928_),
    .B(_2790_),
    .Y(_2929_));
 sky130_fd_sc_hd__nand2_1 _3389_ (.A(_2926_),
    .B(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__a221oi_1 _3390_ (.A1(_2920_),
    .A2(_2921_),
    .B1(_2923_),
    .B2(_2798_),
    .C1(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__clkbuf_8 _3391_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .X(_2932_));
 sky130_fd_sc_hd__inv_2 _3392_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_2933_));
 sky130_fd_sc_hd__or3_1 _3393_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .B(_2754_),
    .C(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__inv_2 _3394_ (.A(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__clkbuf_4 _3395_ (.A(_2935_),
    .X(_2936_));
 sky130_fd_sc_hd__and2_1 _3396_ (.A(_2874_),
    .B(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__buf_1 _3397_ (.A(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__buf_4 _3398_ (.A(_2938_),
    .X(_2939_));
 sky130_fd_sc_hd__and2_1 _3399_ (.A(net36),
    .B(_2860_),
    .X(_2940_));
 sky130_fd_sc_hd__clkbuf_4 _3400_ (.A(_2940_),
    .X(_2941_));
 sky130_fd_sc_hd__nor2_4 _3401_ (.A(_2873_),
    .B(_2876_),
    .Y(_2942_));
 sky130_fd_sc_hd__and2_1 _3402_ (.A(_2942_),
    .B(_2852_),
    .X(_2943_));
 sky130_fd_sc_hd__clkbuf_4 _3403_ (.A(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__nand2_1 _3404_ (.A(_2944_),
    .B(_2788_),
    .Y(_2945_));
 sky130_fd_sc_hd__nor2_4 _3405_ (.A(_2841_),
    .B(_2876_),
    .Y(_2946_));
 sky130_fd_sc_hd__and2_1 _3406_ (.A(_2946_),
    .B(_2852_),
    .X(_2947_));
 sky130_fd_sc_hd__clkbuf_4 _3407_ (.A(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__nand2_1 _3408_ (.A(_2948_),
    .B(_2804_),
    .Y(_2949_));
 sky130_fd_sc_hd__nand2_1 _3409_ (.A(_2945_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__a221oi_1 _3410_ (.A1(_2932_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2794_),
    .C1(_2950_),
    .Y(_2951_));
 sky130_fd_sc_hd__buf_4 _3411_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .X(_2952_));
 sky130_fd_sc_hd__and2_1 _3412_ (.A(_2942_),
    .B(_2835_),
    .X(_2953_));
 sky130_fd_sc_hd__buf_1 _3413_ (.A(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__clkbuf_4 _3414_ (.A(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__clkbuf_8 _3415_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_2956_));
 sky130_fd_sc_hd__and2_1 _3416_ (.A(_2859_),
    .B(_2836_),
    .X(_2957_));
 sky130_fd_sc_hd__clkbuf_2 _3417_ (.A(_2957_),
    .X(_2958_));
 sky130_fd_sc_hd__buf_4 _3418_ (.A(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__and2_1 _3419_ (.A(_2914_),
    .B(_2843_),
    .X(_2960_));
 sky130_fd_sc_hd__clkbuf_4 _3420_ (.A(_2960_),
    .X(_2961_));
 sky130_fd_sc_hd__buf_4 _3421_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .X(_2962_));
 sky130_fd_sc_hd__nand2_1 _3422_ (.A(_2961_),
    .B(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__and2_1 _3423_ (.A(_2946_),
    .B(_2843_),
    .X(_2964_));
 sky130_fd_sc_hd__clkbuf_4 _3424_ (.A(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__clkbuf_8 _3425_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .X(_2966_));
 sky130_fd_sc_hd__nand2_1 _3426_ (.A(_2965_),
    .B(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__nand2_1 _3427_ (.A(_2963_),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__a221oi_1 _3428_ (.A1(_2952_),
    .A2(_2955_),
    .B1(_2956_),
    .B2(_2959_),
    .C1(_2968_),
    .Y(_2969_));
 sky130_fd_sc_hd__and4_1 _3429_ (.A(_2918_),
    .B(_2931_),
    .C(_2951_),
    .D(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__clkbuf_8 _3430_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .X(_2971_));
 sky130_fd_sc_hd__and3_4 _3431_ (.A(_2754_),
    .B(_2822_),
    .C(_2933_),
    .X(_2972_));
 sky130_fd_sc_hd__buf_4 _3432_ (.A(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__and2_1 _3433_ (.A(_2850_),
    .B(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__buf_1 _3434_ (.A(_2974_),
    .X(_2975_));
 sky130_fd_sc_hd__clkbuf_4 _3435_ (.A(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__buf_4 _3436_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .X(_2977_));
 sky130_fd_sc_hd__nor2_4 _3437_ (.A(_2873_),
    .B(_2820_),
    .Y(_2978_));
 sky130_fd_sc_hd__and2_1 _3438_ (.A(_2978_),
    .B(_2836_),
    .X(_2979_));
 sky130_fd_sc_hd__buf_1 _3439_ (.A(_2979_),
    .X(_2980_));
 sky130_fd_sc_hd__clkbuf_4 _3440_ (.A(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__inv_2 _3441_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _3442_ (.A(net36),
    .B(_2973_),
    .Y(_2983_));
 sky130_fd_sc_hd__clkbuf_4 _3443_ (.A(_2983_),
    .X(_2984_));
 sky130_fd_sc_hd__and2_1 _3444_ (.A(_2883_),
    .B(_2836_),
    .X(_2985_));
 sky130_fd_sc_hd__clkbuf_4 _3445_ (.A(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__clkbuf_8 _3446_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .X(_2987_));
 sky130_fd_sc_hd__nand2_1 _3447_ (.A(_2986_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__o21ai_1 _3448_ (.A1(_2982_),
    .A2(_2984_),
    .B1(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__a221oi_1 _3449_ (.A1(_2971_),
    .A2(_2976_),
    .B1(_2977_),
    .B2(_2981_),
    .C1(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__inv_2 _3450_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_2991_));
 sky130_fd_sc_hd__nand2_1 _3451_ (.A(net37),
    .B(_2973_),
    .Y(_2992_));
 sky130_fd_sc_hd__clkbuf_4 _3452_ (.A(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__nand2_1 _3453_ (.A(_2914_),
    .B(_2972_),
    .Y(_2994_));
 sky130_fd_sc_hd__or2b_1 _3454_ (.A(_2994_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_2995_));
 sky130_fd_sc_hd__and2_1 _3455_ (.A(net35),
    .B(_2973_),
    .X(_2996_));
 sky130_fd_sc_hd__clkbuf_4 _3456_ (.A(_2996_),
    .X(_2997_));
 sky130_fd_sc_hd__clkbuf_8 _3457_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_2998_));
 sky130_fd_sc_hd__nand2_1 _3458_ (.A(_2997_),
    .B(_2998_),
    .Y(_2999_));
 sky130_fd_sc_hd__and2_1 _3459_ (.A(_2877_),
    .B(_2936_),
    .X(_3000_));
 sky130_fd_sc_hd__clkbuf_4 _3460_ (.A(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__buf_4 _3461_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .X(_3002_));
 sky130_fd_sc_hd__nand2_1 _3462_ (.A(_3001_),
    .B(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__o2111a_1 _3463_ (.A1(_2991_),
    .A2(_2993_),
    .B1(_2995_),
    .C1(_2999_),
    .D1(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__buf_4 _3464_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .X(_3005_));
 sky130_fd_sc_hd__and2_1 _3465_ (.A(_2946_),
    .B(_2835_),
    .X(_3006_));
 sky130_fd_sc_hd__buf_1 _3466_ (.A(_3006_),
    .X(_3007_));
 sky130_fd_sc_hd__buf_4 _3467_ (.A(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__buf_4 _3468_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .X(_3009_));
 sky130_fd_sc_hd__and2_1 _3469_ (.A(_2855_),
    .B(_2835_),
    .X(_3010_));
 sky130_fd_sc_hd__buf_1 _3470_ (.A(_3010_),
    .X(_3011_));
 sky130_fd_sc_hd__buf_4 _3471_ (.A(_3011_),
    .X(_3012_));
 sky130_fd_sc_hd__buf_4 _3472_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_3013_));
 sky130_fd_sc_hd__inv_2 _3473_ (.A(_3013_),
    .Y(_3014_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(_2850_),
    .B(_2836_),
    .Y(_3015_));
 sky130_fd_sc_hd__clkbuf_4 _3475_ (.A(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__clkbuf_8 _3476_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_3017_));
 sky130_fd_sc_hd__inv_2 _3477_ (.A(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__and3_2 _3478_ (.A(_2754_),
    .B(_2933_),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3019_));
 sky130_fd_sc_hd__clkbuf_4 _3479_ (.A(_3019_),
    .X(_3020_));
 sky130_fd_sc_hd__nand2_1 _3480_ (.A(_2978_),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__clkbuf_4 _3481_ (.A(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__o22ai_1 _3482_ (.A1(_3014_),
    .A2(_3016_),
    .B1(_3018_),
    .B2(_3022_),
    .Y(_3023_));
 sky130_fd_sc_hd__a221oi_1 _3483_ (.A1(_3005_),
    .A2(_3008_),
    .B1(_3009_),
    .B2(_3012_),
    .C1(_3023_),
    .Y(_3024_));
 sky130_fd_sc_hd__and3_2 _3484_ (.A(_2822_),
    .B(_2933_),
    .C(\egd_top.BitStream_buffer.pc[6] ),
    .X(_3025_));
 sky130_fd_sc_hd__clkbuf_4 _3485_ (.A(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__and2_1 _3486_ (.A(_2855_),
    .B(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__clkbuf_4 _3487_ (.A(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__clkbuf_8 _3488_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_3029_));
 sky130_fd_sc_hd__clkbuf_8 _3489_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_3030_));
 sky130_fd_sc_hd__and2_1 _3490_ (.A(_2859_),
    .B(_3026_),
    .X(_3031_));
 sky130_fd_sc_hd__buf_1 _3491_ (.A(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__buf_4 _3492_ (.A(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__and2_1 _3493_ (.A(_2753_),
    .B(_2936_),
    .X(_3034_));
 sky130_fd_sc_hd__clkbuf_4 _3494_ (.A(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__clkbuf_8 _3495_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .X(_3036_));
 sky130_fd_sc_hd__nand2_1 _3496_ (.A(_3035_),
    .B(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__and2_1 _3497_ (.A(_2946_),
    .B(_3026_),
    .X(_3038_));
 sky130_fd_sc_hd__clkbuf_4 _3498_ (.A(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__nand2_1 _3499_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_3040_));
 sky130_fd_sc_hd__nand2_1 _3500_ (.A(_3037_),
    .B(_3040_),
    .Y(_3041_));
 sky130_fd_sc_hd__a221oi_1 _3501_ (.A1(_3028_),
    .A2(_3029_),
    .B1(_3030_),
    .B2(_3033_),
    .C1(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__and4_1 _3502_ (.A(_2990_),
    .B(_3004_),
    .C(_3024_),
    .D(_3042_),
    .X(_3043_));
 sky130_fd_sc_hd__buf_4 _3503_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .X(_3044_));
 sky130_fd_sc_hd__and2_1 _3504_ (.A(_2978_),
    .B(_2755_),
    .X(_3045_));
 sky130_fd_sc_hd__clkbuf_2 _3505_ (.A(_3045_),
    .X(_3046_));
 sky130_fd_sc_hd__buf_4 _3506_ (.A(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__and2_2 _3507_ (.A(net38),
    .B(_3020_),
    .X(_3048_));
 sky130_fd_sc_hd__buf_4 _3508_ (.A(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__buf_4 _3509_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_3050_));
 sky130_fd_sc_hd__and2_1 _3510_ (.A(_2753_),
    .B(_3019_),
    .X(_3051_));
 sky130_fd_sc_hd__clkbuf_4 _3511_ (.A(_3051_),
    .X(_3052_));
 sky130_fd_sc_hd__buf_4 _3512_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_3053_));
 sky130_fd_sc_hd__nand2_1 _3513_ (.A(_3052_),
    .B(_3053_),
    .Y(_3054_));
 sky130_fd_sc_hd__buf_2 _3514_ (.A(_2755_),
    .X(_3055_));
 sky130_fd_sc_hd__and2_1 _3515_ (.A(_2874_),
    .B(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__buf_4 _3516_ (.A(_3056_),
    .X(_3057_));
 sky130_fd_sc_hd__buf_4 _3517_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_3058_));
 sky130_fd_sc_hd__nand2_1 _3518_ (.A(_3057_),
    .B(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__nand2_1 _3519_ (.A(_3054_),
    .B(_3059_),
    .Y(_3060_));
 sky130_fd_sc_hd__a221oi_1 _3520_ (.A1(_3044_),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_3050_),
    .C1(_3060_),
    .Y(_3061_));
 sky130_fd_sc_hd__and2_1 _3521_ (.A(_2753_),
    .B(_3026_),
    .X(_3062_));
 sky130_fd_sc_hd__clkbuf_4 _3522_ (.A(_3062_),
    .X(_3063_));
 sky130_fd_sc_hd__clkbuf_8 _3523_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_3064_));
 sky130_fd_sc_hd__and2_1 _3524_ (.A(net38),
    .B(_3026_),
    .X(_3065_));
 sky130_fd_sc_hd__clkbuf_4 _3525_ (.A(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__clkbuf_8 _3526_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .X(_3067_));
 sky130_fd_sc_hd__and2_1 _3527_ (.A(_2883_),
    .B(_2852_),
    .X(_3068_));
 sky130_fd_sc_hd__clkbuf_4 _3528_ (.A(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__nand2_1 _3529_ (.A(_3069_),
    .B(_2802_),
    .Y(_3070_));
 sky130_fd_sc_hd__and2_1 _3530_ (.A(_2842_),
    .B(_3026_),
    .X(_3071_));
 sky130_fd_sc_hd__clkbuf_4 _3531_ (.A(_3071_),
    .X(_3072_));
 sky130_fd_sc_hd__nand2_1 _3532_ (.A(_3072_),
    .B(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_3073_));
 sky130_fd_sc_hd__nand2_1 _3533_ (.A(_3070_),
    .B(_3073_),
    .Y(_3074_));
 sky130_fd_sc_hd__a221oi_1 _3534_ (.A1(_3063_),
    .A2(_3064_),
    .B1(_3066_),
    .B2(_3067_),
    .C1(_3074_),
    .Y(_3075_));
 sky130_fd_sc_hd__and2_1 _3535_ (.A(_2874_),
    .B(_2973_),
    .X(_3076_));
 sky130_fd_sc_hd__clkbuf_4 _3536_ (.A(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__clkbuf_8 _3537_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_3078_));
 sky130_fd_sc_hd__buf_4 _3538_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .X(_3079_));
 sky130_fd_sc_hd__and2_1 _3539_ (.A(_2859_),
    .B(_2755_),
    .X(_3080_));
 sky130_fd_sc_hd__clkbuf_2 _3540_ (.A(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__buf_4 _3541_ (.A(_3081_),
    .X(_3082_));
 sky130_fd_sc_hd__clkbuf_8 _3542_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .X(_3083_));
 sky130_fd_sc_hd__inv_2 _3543_ (.A(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__nand2_1 _3544_ (.A(_2859_),
    .B(_2973_),
    .Y(_3085_));
 sky130_fd_sc_hd__clkbuf_4 _3545_ (.A(_3085_),
    .X(_3086_));
 sky130_fd_sc_hd__and2_1 _3546_ (.A(_2942_),
    .B(_2973_),
    .X(_3087_));
 sky130_fd_sc_hd__clkbuf_4 _3547_ (.A(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__nand2_1 _3548_ (.A(_3088_),
    .B(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .Y(_3089_));
 sky130_fd_sc_hd__o21ai_1 _3549_ (.A1(_3084_),
    .A2(_3086_),
    .B1(_3089_),
    .Y(_3090_));
 sky130_fd_sc_hd__a221oi_1 _3550_ (.A1(_3077_),
    .A2(_3078_),
    .B1(_3079_),
    .B2(_3082_),
    .C1(_3090_),
    .Y(_3091_));
 sky130_fd_sc_hd__clkbuf_8 _3551_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_3092_));
 sky130_fd_sc_hd__and2_1 _3552_ (.A(_2842_),
    .B(_3019_),
    .X(_3093_));
 sky130_fd_sc_hd__buf_1 _3553_ (.A(_3093_),
    .X(_3094_));
 sky130_fd_sc_hd__clkbuf_4 _3554_ (.A(_3094_),
    .X(_3095_));
 sky130_fd_sc_hd__and2_1 _3555_ (.A(net38),
    .B(_2936_),
    .X(_3096_));
 sky130_fd_sc_hd__clkbuf_4 _3556_ (.A(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__clkbuf_8 _3557_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .X(_3098_));
 sky130_fd_sc_hd__and2_1 _3558_ (.A(_2877_),
    .B(_3026_),
    .X(_3099_));
 sky130_fd_sc_hd__clkbuf_4 _3559_ (.A(_3099_),
    .X(_3100_));
 sky130_fd_sc_hd__nand2_1 _3560_ (.A(_3100_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_3101_));
 sky130_fd_sc_hd__and2_1 _3561_ (.A(_2842_),
    .B(_2936_),
    .X(_3102_));
 sky130_fd_sc_hd__clkbuf_4 _3562_ (.A(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__clkbuf_8 _3563_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_3104_));
 sky130_fd_sc_hd__nand2_1 _3564_ (.A(_3103_),
    .B(_3104_),
    .Y(_3105_));
 sky130_fd_sc_hd__nand2_1 _3565_ (.A(_3101_),
    .B(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__a221oi_1 _3566_ (.A1(_3092_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_3098_),
    .C1(_3106_),
    .Y(_3107_));
 sky130_fd_sc_hd__and4_1 _3567_ (.A(_3061_),
    .B(_3075_),
    .C(_3091_),
    .D(_3107_),
    .X(_3108_));
 sky130_fd_sc_hd__and4_1 _3568_ (.A(_2898_),
    .B(_2970_),
    .C(_3043_),
    .D(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__o41a_1 _3569_ (.A1(\egd_top.BitStream_buffer.pc[2] ),
    .A2(\egd_top.BitStream_buffer.pc[3] ),
    .A3(\egd_top.BitStream_buffer.pc[1] ),
    .A4(\egd_top.BitStream_buffer.pc[0] ),
    .B1(_2973_),
    .X(_3110_));
 sky130_fd_sc_hd__or4_1 _3570_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .D(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__clkbuf_4 _3571_ (.A(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__buf_4 _3572_ (.A(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__buf_4 _3573_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_3114_));
 sky130_fd_sc_hd__and2_1 _3574_ (.A(_2914_),
    .B(_3055_),
    .X(_3115_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3575_ (.A(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__buf_4 _3576_ (.A(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__buf_4 _3577_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .X(_3118_));
 sky130_fd_sc_hd__and2_1 _3578_ (.A(_2946_),
    .B(_3055_),
    .X(_3119_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3579_ (.A(_3119_),
    .X(_3120_));
 sky130_fd_sc_hd__buf_4 _3580_ (.A(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__inv_2 _3581_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_3122_));
 sky130_fd_sc_hd__nand2_1 _3582_ (.A(_2829_),
    .B(_3055_),
    .Y(_3123_));
 sky130_fd_sc_hd__clkbuf_4 _3583_ (.A(_3123_),
    .X(_3124_));
 sky130_fd_sc_hd__and2_1 _3584_ (.A(net38),
    .B(_3055_),
    .X(_3125_));
 sky130_fd_sc_hd__clkbuf_4 _3585_ (.A(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__buf_4 _3586_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_3127_));
 sky130_fd_sc_hd__nand2_1 _3587_ (.A(_3126_),
    .B(_3127_),
    .Y(_3128_));
 sky130_fd_sc_hd__o21ai_1 _3588_ (.A1(_3122_),
    .A2(_3124_),
    .B1(_3128_),
    .Y(_3129_));
 sky130_fd_sc_hd__a221oi_2 _3589_ (.A1(_3114_),
    .A2(_3117_),
    .B1(_3118_),
    .B2(_3121_),
    .C1(_3129_),
    .Y(_3130_));
 sky130_fd_sc_hd__inv_2 _3590_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_3131_));
 sky130_fd_sc_hd__nand2_1 _3591_ (.A(_2834_),
    .B(_3055_),
    .Y(_3132_));
 sky130_fd_sc_hd__clkbuf_4 _3592_ (.A(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__buf_6 _3593_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .X(_3134_));
 sky130_fd_sc_hd__inv_2 _3594_ (.A(_3134_),
    .Y(_3135_));
 sky130_fd_sc_hd__nand2_1 _3595_ (.A(_2855_),
    .B(_2972_),
    .Y(_3136_));
 sky130_fd_sc_hd__buf_2 _3596_ (.A(_3136_),
    .X(_3137_));
 sky130_fd_sc_hd__or2_1 _3597_ (.A(_3135_),
    .B(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__inv_2 _3598_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_3139_));
 sky130_fd_sc_hd__nand2_1 _3599_ (.A(_2883_),
    .B(_2972_),
    .Y(_3140_));
 sky130_fd_sc_hd__buf_2 _3600_ (.A(_3140_),
    .X(_3141_));
 sky130_fd_sc_hd__or2_1 _3601_ (.A(_3139_),
    .B(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__and2_1 _3602_ (.A(_2900_),
    .B(_3055_),
    .X(_3143_));
 sky130_fd_sc_hd__clkbuf_4 _3603_ (.A(_3143_),
    .X(_3144_));
 sky130_fd_sc_hd__nand2_1 _3604_ (.A(_3144_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_3145_));
 sky130_fd_sc_hd__o2111a_1 _3605_ (.A1(_3131_),
    .A2(_3133_),
    .B1(_3138_),
    .C1(_3142_),
    .D1(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__buf_4 _3606_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_3147_));
 sky130_fd_sc_hd__and2_1 _3607_ (.A(_2877_),
    .B(_2835_),
    .X(_3148_));
 sky130_fd_sc_hd__clkbuf_2 _3608_ (.A(_3148_),
    .X(_3149_));
 sky130_fd_sc_hd__clkbuf_4 _3609_ (.A(_3149_),
    .X(_3150_));
 sky130_fd_sc_hd__and2_2 _3610_ (.A(net37),
    .B(_3026_),
    .X(_3151_));
 sky130_fd_sc_hd__clkbuf_4 _3611_ (.A(_3151_),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_8 _3612_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _3613_ (.A(_2753_),
    .B(_2836_),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_4 _3614_ (.A(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__buf_4 _3615_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _3616_ (.A(_0325_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__and2_1 _3617_ (.A(_2946_),
    .B(_2973_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _3618_ (.A(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_8 _3619_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _3620_ (.A(_0329_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2_1 _3621_ (.A(_0327_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__a221oi_1 _3622_ (.A1(_3147_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0323_),
    .C1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__buf_4 _3623_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_0334_));
 sky130_fd_sc_hd__and2_1 _3624_ (.A(_2942_),
    .B(_3019_),
    .X(_0335_));
 sky130_fd_sc_hd__buf_1 _3625_ (.A(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_4 _3626_ (.A(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_8 _3627_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _3628_ (.A(_2874_),
    .B(_3019_),
    .X(_0339_));
 sky130_fd_sc_hd__buf_1 _3629_ (.A(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_4 _3630_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__inv_2 _3631_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _3632_ (.A(_2842_),
    .B(_3055_),
    .Y(_0343_));
 sky130_fd_sc_hd__clkbuf_4 _3633_ (.A(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_8 _3634_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_0345_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand2_1 _3636_ (.A(_2859_),
    .B(_3020_),
    .Y(_0347_));
 sky130_fd_sc_hd__clkbuf_4 _3637_ (.A(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__o22ai_1 _3638_ (.A1(_0342_),
    .A2(_0344_),
    .B1(_0346_),
    .B2(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__a221oi_1 _3639_ (.A1(_0334_),
    .A2(_0337_),
    .B1(_0338_),
    .B2(_0341_),
    .C1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__and4_1 _3640_ (.A(_3130_),
    .B(_3146_),
    .C(_0333_),
    .D(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_8 _3641_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_0352_));
 sky130_fd_sc_hd__and2_1 _3642_ (.A(_2883_),
    .B(_3025_),
    .X(_0353_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3643_ (.A(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__buf_4 _3644_ (.A(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _3645_ (.A(_2834_),
    .B(_3020_),
    .X(_0356_));
 sky130_fd_sc_hd__buf_4 _3646_ (.A(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_8 _3647_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _3648_ (.A(_2883_),
    .B(_3055_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_4 _3649_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__nand2_1 _3650_ (.A(_0360_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0361_));
 sky130_fd_sc_hd__and2_1 _3651_ (.A(_2855_),
    .B(_3055_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_4 _3652_ (.A(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__buf_4 _3653_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _3654_ (.A(_0363_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_1 _3655_ (.A(_0361_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__a221oi_2 _3656_ (.A1(_0352_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0358_),
    .C1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_1 _3657_ (.A(_2834_),
    .B(_2935_),
    .Y(_0368_));
 sky130_fd_sc_hd__clkbuf_4 _3658_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__or2b_1 _3659_ (.A(_0369_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_0370_));
 sky130_fd_sc_hd__and2_1 _3660_ (.A(_2942_),
    .B(_2936_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_4 _3661_ (.A(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__nand2_1 _3662_ (.A(_0372_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0373_));
 sky130_fd_sc_hd__and2_1 _3663_ (.A(_2914_),
    .B(_2935_),
    .X(_0374_));
 sky130_fd_sc_hd__buf_4 _3664_ (.A(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__nand2_1 _3665_ (.A(_0375_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0376_));
 sky130_fd_sc_hd__and2_1 _3666_ (.A(_2883_),
    .B(_2935_),
    .X(_0377_));
 sky130_fd_sc_hd__buf_4 _3667_ (.A(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__buf_4 _3668_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _3669_ (.A(_0378_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__and4_1 _3670_ (.A(_0370_),
    .B(_0373_),
    .C(_0376_),
    .D(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _3671_ (.A(_2914_),
    .B(_3020_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_4 _3672_ (.A(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_8 _3673_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_0384_));
 sky130_fd_sc_hd__buf_4 _3674_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _3675_ (.A(_2874_),
    .B(_3025_),
    .X(_0386_));
 sky130_fd_sc_hd__buf_1 _3676_ (.A(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_4 _3677_ (.A(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _3678_ (.A(_2850_),
    .B(_2755_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_4 _3679_ (.A(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__buf_4 _3680_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .X(_0391_));
 sky130_fd_sc_hd__nand2_1 _3681_ (.A(_0390_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__and2_1 _3682_ (.A(_2877_),
    .B(_2755_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_4 _3683_ (.A(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__buf_4 _3684_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _3685_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__nand2_1 _3686_ (.A(_0392_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__a221oi_1 _3687_ (.A1(_0383_),
    .A2(_0384_),
    .B1(_0385_),
    .B2(_0388_),
    .C1(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(_2942_),
    .B(_3025_),
    .Y(_0399_));
 sky130_fd_sc_hd__inv_2 _3689_ (.A(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__clkbuf_4 _3690_ (.A(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__nand2_1 _3691_ (.A(_2834_),
    .B(_3025_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _3692_ (.A(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__clkbuf_4 _3693_ (.A(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__a22o_1 _3694_ (.A1(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _3695_ (.A(_2900_),
    .B(_2935_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_4 _3696_ (.A(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _3697_ (.A(_2829_),
    .B(_2936_),
    .X(_0408_));
 sky130_fd_sc_hd__buf_4 _3698_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_8 _3699_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0410_));
 sky130_fd_sc_hd__a22o_1 _3700_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .B1(_0409_),
    .B2(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _3701_ (.A(_0405_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__and4_1 _3702_ (.A(_0367_),
    .B(_0381_),
    .C(_0398_),
    .D(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _3703_ (.A(_2914_),
    .B(_3026_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_4 _3704_ (.A(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__buf_4 _3705_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _3706_ (.A(net35),
    .B(_3026_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_4 _3707_ (.A(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__buf_4 _3708_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_0419_));
 sky130_fd_sc_hd__and2_1 _3709_ (.A(_2850_),
    .B(_3026_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_4 _3710_ (.A(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_8 _3711_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _3712_ (.A(_0421_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__and2_1 _3713_ (.A(_2978_),
    .B(_2936_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_4 _3714_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_8 _3715_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_0426_));
 sky130_fd_sc_hd__nand2_1 _3716_ (.A(_0425_),
    .B(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__nand2_1 _3717_ (.A(_0423_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__a221oi_1 _3718_ (.A1(_0415_),
    .A2(_0416_),
    .B1(_0418_),
    .B2(_0419_),
    .C1(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__clkbuf_8 _3719_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .X(_0430_));
 sky130_fd_sc_hd__and2_1 _3720_ (.A(_2842_),
    .B(_2972_),
    .X(_0431_));
 sky130_fd_sc_hd__buf_1 _3721_ (.A(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_4 _3722_ (.A(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _3723_ (.A(net38),
    .B(_2973_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_4 _3724_ (.A(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__buf_4 _3725_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_0436_));
 sky130_fd_sc_hd__and2_1 _3726_ (.A(_2850_),
    .B(_2936_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_4 _3727_ (.A(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__buf_4 _3728_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_1 _3729_ (.A(_0438_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__and2_1 _3730_ (.A(_2978_),
    .B(_2824_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_4 _3731_ (.A(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__buf_4 _3732_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_1 _3733_ (.A(_0442_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _3734_ (.A(_0440_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__a221oi_1 _3735_ (.A1(_0430_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_0436_),
    .C1(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__clkbuf_8 _3736_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .X(_0447_));
 sky130_fd_sc_hd__inv_2 _3737_ (.A(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _3738_ (.A(_2842_),
    .B(_2836_),
    .Y(_0449_));
 sky130_fd_sc_hd__clkbuf_4 _3739_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_4 _3740_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .X(_0451_));
 sky130_fd_sc_hd__inv_2 _3741_ (.A(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand2_1 _3742_ (.A(_2821_),
    .B(_2836_),
    .Y(_0453_));
 sky130_fd_sc_hd__clkbuf_4 _3743_ (.A(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__o22ai_1 _3744_ (.A1(_0448_),
    .A2(_0450_),
    .B1(_0452_),
    .B2(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__and2_1 _3745_ (.A(_2877_),
    .B(_2973_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_8 _3746_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .X(_0457_));
 sky130_fd_sc_hd__and2_1 _3747_ (.A(_2753_),
    .B(_2973_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_8 _3748_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _3749_ (.A1(_0456_),
    .A2(_0457_),
    .B1(_0458_),
    .B2(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_1 _3750_ (.A(_0455_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_2 _3751_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _3752_ (.A(_2942_),
    .B(_2843_),
    .Y(_0463_));
 sky130_fd_sc_hd__clkbuf_4 _3753_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__inv_2 _3754_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_1 _3755_ (.A(_2859_),
    .B(_2936_),
    .Y(_0466_));
 sky130_fd_sc_hd__clkbuf_4 _3756_ (.A(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__o22ai_1 _3757_ (.A1(_0462_),
    .A2(_0464_),
    .B1(_0465_),
    .B2(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__and2_1 _3758_ (.A(_2946_),
    .B(_2936_),
    .X(_0469_));
 sky130_fd_sc_hd__and2_1 _3759_ (.A(_2855_),
    .B(_2936_),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_8 _3760_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _3761_ (.A1(_0469_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .B1(_0470_),
    .B2(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__nor2_1 _3762_ (.A(_0468_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__and4_1 _3763_ (.A(_0429_),
    .B(_0446_),
    .C(_0461_),
    .D(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__buf_4 _3764_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _3765_ (.A(_2978_),
    .B(_3026_),
    .X(_0476_));
 sky130_fd_sc_hd__buf_1 _3766_ (.A(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_4 _3767_ (.A(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_4 _3768_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .X(_0479_));
 sky130_fd_sc_hd__buf_4 _3769_ (.A(_2757_),
    .X(_0480_));
 sky130_fd_sc_hd__inv_2 _3770_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_0481_));
 sky130_fd_sc_hd__nand2_1 _3771_ (.A(_2946_),
    .B(_3020_),
    .Y(_0482_));
 sky130_fd_sc_hd__clkbuf_4 _3772_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__buf_4 _3773_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_0484_));
 sky130_fd_sc_hd__inv_2 _3774_ (.A(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__nand2_1 _3775_ (.A(_2850_),
    .B(_3020_),
    .Y(_0486_));
 sky130_fd_sc_hd__clkbuf_4 _3776_ (.A(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__o22ai_1 _3777_ (.A1(_0481_),
    .A2(_0483_),
    .B1(_0485_),
    .B2(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__a221oi_2 _3778_ (.A1(_0475_),
    .A2(_0478_),
    .B1(_0479_),
    .B2(_0480_),
    .C1(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _3779_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _3780_ (.A(_2883_),
    .B(_3020_),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_2 _3781_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_0492_));
 sky130_fd_sc_hd__nand2_1 _3782_ (.A(_2855_),
    .B(_3020_),
    .Y(_0493_));
 sky130_fd_sc_hd__o22ai_1 _3783_ (.A1(_0490_),
    .A2(_0491_),
    .B1(_0492_),
    .B2(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__and2_1 _3784_ (.A(net35),
    .B(_3020_),
    .X(_0495_));
 sky130_fd_sc_hd__and2_1 _3785_ (.A(net37),
    .B(_3020_),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _3786_ (.A1(_0495_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .B1(_0496_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_1 _3787_ (.A(_0494_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _3788_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _3789_ (.A(_2874_),
    .B(_2843_),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _3790_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_0501_));
 sky130_fd_sc_hd__nand2_2 _3791_ (.A(_2859_),
    .B(_2843_),
    .Y(_0502_));
 sky130_fd_sc_hd__clkbuf_4 _3792_ (.A(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o22ai_1 _3793_ (.A1(_0499_),
    .A2(_0500_),
    .B1(_0501_),
    .B2(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__and2_1 _3794_ (.A(_2978_),
    .B(_2852_),
    .X(_0505_));
 sky130_fd_sc_hd__and2_1 _3795_ (.A(_2753_),
    .B(_2824_),
    .X(_0506_));
 sky130_fd_sc_hd__buf_4 _3796_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .X(_0507_));
 sky130_fd_sc_hd__a22o_1 _3797_ (.A1(_0505_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .B1(_0506_),
    .B2(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__nor2_1 _3798_ (.A(_0504_),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__buf_4 _3799_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_0510_));
 sky130_fd_sc_hd__inv_2 _3800_ (.A(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _3801_ (.A(_2877_),
    .B(_3020_),
    .Y(_0512_));
 sky130_fd_sc_hd__buf_4 _3802_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_0513_));
 sky130_fd_sc_hd__inv_2 _3803_ (.A(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_1 _3804_ (.A(_2942_),
    .B(_3055_),
    .Y(_0515_));
 sky130_fd_sc_hd__o22ai_1 _3805_ (.A1(_0511_),
    .A2(_0512_),
    .B1(_0514_),
    .B2(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__and2_1 _3806_ (.A(_2877_),
    .B(_2852_),
    .X(_0517_));
 sky130_fd_sc_hd__and2_1 _3807_ (.A(_2753_),
    .B(_2852_),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _3808_ (.A1(_0517_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .B1(_0518_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_0519_));
 sky130_fd_sc_hd__nor2_1 _3809_ (.A(_0516_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__and4_1 _3810_ (.A(_0489_),
    .B(_0498_),
    .C(_0509_),
    .D(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__and4_1 _3811_ (.A(_0351_),
    .B(_0413_),
    .C(_0474_),
    .D(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__nand3_2 _3812_ (.A(_3109_),
    .B(_3113_),
    .C(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__buf_4 _3813_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_4 _3814_ (.A(_3112_),
    .X(_0525_));
 sky130_fd_sc_hd__o21a_1 _3815_ (.A1(_0524_),
    .A2(_0525_),
    .B1(_2776_),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _3816_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B1(_0523_),
    .B2(_0526_),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_1 _3817_ (.A(_2838_),
    .B(_2899_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _3818_ (.A(_2845_),
    .B(_2886_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_1 _3819_ (.A(_0527_),
    .B(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__a221oi_2 _3820_ (.A1(_2865_),
    .A2(_2827_),
    .B1(_2846_),
    .B2(_2832_),
    .C1(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__a22o_1 _3821_ (.A1(_2854_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .B1(_2857_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _3822_ (.A1(_2812_),
    .A2(_2862_),
    .B1(_2864_),
    .B2(_2921_),
    .X(_0532_));
 sky130_fd_sc_hd__nor2_1 _3823_ (.A(_0531_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _3824_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _3825_ (.A(_2879_),
    .B(_0507_),
    .Y(_0535_));
 sky130_fd_sc_hd__o221a_1 _3826_ (.A1(_0501_),
    .A2(_2870_),
    .B1(_0534_),
    .B2(_2875_),
    .C1(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_8 _3827_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .X(_0537_));
 sky130_fd_sc_hd__nand2_1 _3828_ (.A(_2890_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _3829_ (.A(_2894_),
    .B(_2802_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _3830_ (.A(_0538_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__a221oi_1 _3831_ (.A1(_2885_),
    .A2(_2966_),
    .B1(_2888_),
    .B2(_2794_),
    .C1(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__and4_1 _3832_ (.A(_0530_),
    .B(_0533_),
    .C(_0536_),
    .D(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__inv_2 _3833_ (.A(_2952_),
    .Y(_0543_));
 sky130_fd_sc_hd__o22ai_1 _3834_ (.A1(_0543_),
    .A2(_2911_),
    .B1(_0452_),
    .B2(_2916_),
    .Y(_0544_));
 sky130_fd_sc_hd__a221oi_1 _3835_ (.A1(_2904_),
    .A2(_2903_),
    .B1(_0447_),
    .B2(_2907_),
    .C1(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _3836_ (.A(_2925_),
    .B(_2798_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _3837_ (.A(_2928_),
    .B(_2792_),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _3838_ (.A(_0546_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a221oi_1 _3839_ (.A1(_2920_),
    .A2(_2828_),
    .B1(_2923_),
    .B2(_2800_),
    .C1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__clkbuf_8 _3840_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_1 _3841_ (.A(_2944_),
    .B(_2790_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _3842_ (.A(_2948_),
    .B(_2806_),
    .Y(_0552_));
 sky130_fd_sc_hd__nand2_1 _3843_ (.A(_0551_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__a221oi_1 _3844_ (.A1(_0550_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2796_),
    .C1(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _3845_ (.A(_2961_),
    .B(_2817_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand2_1 _3846_ (.A(_2965_),
    .B(_2891_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _3847_ (.A(_0555_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__a221oi_1 _3848_ (.A1(_2912_),
    .A2(_2955_),
    .B1(_3147_),
    .B2(_2959_),
    .C1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__and4_1 _3849_ (.A(_0545_),
    .B(_0549_),
    .C(_0554_),
    .D(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__inv_2 _3850_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_1 _3851_ (.A(_2986_),
    .B(_3005_),
    .Y(_0561_));
 sky130_fd_sc_hd__o21ai_1 _3852_ (.A1(_0560_),
    .A2(_2984_),
    .B1(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__a221oi_1 _3853_ (.A1(_3083_),
    .A2(_2976_),
    .B1(_2908_),
    .B2(_2981_),
    .C1(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_2 _3854_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0564_));
 sky130_fd_sc_hd__or2b_1 _3855_ (.A(_2994_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_0565_));
 sky130_fd_sc_hd__buf_4 _3856_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .X(_0566_));
 sky130_fd_sc_hd__nand2_1 _3857_ (.A(_2997_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_3001_),
    .B(_3036_),
    .Y(_0568_));
 sky130_fd_sc_hd__o2111a_1 _3859_ (.A1(_0564_),
    .A2(_2993_),
    .B1(_0565_),
    .C1(_0567_),
    .D1(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__inv_2 _3860_ (.A(_2956_),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_2 _3861_ (.A(_0338_),
    .Y(_0571_));
 sky130_fd_sc_hd__o22ai_1 _3862_ (.A1(_0570_),
    .A2(_3016_),
    .B1(_0571_),
    .B2(_3022_),
    .Y(_0572_));
 sky130_fd_sc_hd__a221oi_1 _3863_ (.A1(_3009_),
    .A2(_3008_),
    .B1(_3013_),
    .B2(_3012_),
    .C1(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__clkbuf_8 _3864_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_0574_));
 sky130_fd_sc_hd__nand2_1 _3865_ (.A(_3035_),
    .B(_0443_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _3866_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _3867_ (.A(_0575_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__a221oi_1 _3868_ (.A1(_3028_),
    .A2(_0422_),
    .B1(_0574_),
    .B2(_3033_),
    .C1(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__and4_1 _3869_ (.A(_0563_),
    .B(_0569_),
    .C(_0573_),
    .D(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__nand2_1 _3870_ (.A(_3052_),
    .B(_3044_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_1 _3871_ (.A(_3057_),
    .B(_0513_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _3872_ (.A(_0580_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__a221oi_2 _3873_ (.A1(_3058_),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0358_),
    .C1(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__clkbuf_8 _3874_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_0584_));
 sky130_fd_sc_hd__nand2_1 _3875_ (.A(_3069_),
    .B(_2804_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_1 _3876_ (.A(_3072_),
    .B(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__a221oi_1 _3878_ (.A1(_3063_),
    .A2(_0426_),
    .B1(_3066_),
    .B2(_0584_),
    .C1(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__buf_4 _3879_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_0589_));
 sky130_fd_sc_hd__inv_2 _3880_ (.A(_0457_),
    .Y(_0590_));
 sky130_fd_sc_hd__clkbuf_8 _3881_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_0591_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(_3088_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__o21ai_1 _3883_ (.A1(_0590_),
    .A2(_3086_),
    .B1(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a221oi_1 _3884_ (.A1(_3077_),
    .A2(_0589_),
    .B1(_0395_),
    .B2(_3082_),
    .C1(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__buf_6 _3885_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_8 _3886_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_0596_));
 sky130_fd_sc_hd__nand2_1 _3887_ (.A(_3100_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _3888_ (.A(_3103_),
    .B(_0379_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2_1 _3889_ (.A(_0597_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__a221oi_1 _3890_ (.A1(_0595_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0596_),
    .C1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__and4_2 _3891_ (.A(_0583_),
    .B(_0588_),
    .C(_0594_),
    .D(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__and4_1 _3892_ (.A(_0542_),
    .B(_0559_),
    .C(_0579_),
    .D(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__nand2_1 _3893_ (.A(_3126_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_0603_));
 sky130_fd_sc_hd__o21ai_1 _3894_ (.A1(_0342_),
    .A2(_3124_),
    .B1(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__a221oi_2 _3895_ (.A1(_3127_),
    .A2(_3117_),
    .B1(_0364_),
    .B2(_3121_),
    .C1(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__inv_2 _3896_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0606_));
 sky130_fd_sc_hd__inv_2 _3897_ (.A(_2971_),
    .Y(_0607_));
 sky130_fd_sc_hd__or2_1 _3898_ (.A(_0607_),
    .B(_3137_),
    .X(_0608_));
 sky130_fd_sc_hd__inv_2 _3899_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0609_));
 sky130_fd_sc_hd__or2_1 _3900_ (.A(_0609_),
    .B(_3141_),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_1 _3901_ (.A(_3144_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_0611_));
 sky130_fd_sc_hd__o2111a_1 _3902_ (.A1(_0606_),
    .A2(_3133_),
    .B1(_0608_),
    .C1(_0610_),
    .D1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_8 _3903_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_1 _3904_ (.A(_0325_),
    .B(_3017_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_1 _3905_ (.A(_0329_),
    .B(_3134_),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_1 _3906_ (.A(_0614_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a221oi_1 _3907_ (.A1(_0326_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0613_),
    .C1(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__clkinv_4 _3908_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0618_));
 sky130_fd_sc_hd__o22ai_1 _3909_ (.A1(_0618_),
    .A2(_0344_),
    .B1(_0511_),
    .B2(_0348_),
    .Y(_0619_));
 sky130_fd_sc_hd__a221oi_1 _3910_ (.A1(_0384_),
    .A2(_0337_),
    .B1(_0334_),
    .B2(_0341_),
    .C1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__and4_1 _3911_ (.A(_0605_),
    .B(_0612_),
    .C(_0617_),
    .D(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_8 _3912_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_8 _3913_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_0623_));
 sky130_fd_sc_hd__nand2_1 _3914_ (.A(_0360_),
    .B(_3118_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _3915_ (.A(_0363_),
    .B(_0391_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _3916_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__a221oi_2 _3917_ (.A1(_0622_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0623_),
    .C1(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__or2b_1 _3918_ (.A(_0369_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_0628_));
 sky130_fd_sc_hd__nand2_1 _3919_ (.A(_0372_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _3920_ (.A(_0375_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0630_));
 sky130_fd_sc_hd__clkbuf_8 _3921_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_0631_));
 sky130_fd_sc_hd__nand2_1 _3922_ (.A(_0378_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__and4_1 _3923_ (.A(_0628_),
    .B(_0629_),
    .C(_0630_),
    .D(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__buf_4 _3924_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _3925_ (.A(_0390_),
    .B(_3079_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2_1 _3926_ (.A(_0394_),
    .B(_0479_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_0635_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a221oi_1 _3928_ (.A1(_0383_),
    .A2(_3050_),
    .B1(_0634_),
    .B2(_0388_),
    .C1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__a22o_1 _3929_ (.A1(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _3930_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .B1(_0409_),
    .B2(_3104_),
    .X(_0640_));
 sky130_fd_sc_hd__nor2_1 _3931_ (.A(_0639_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__and4_1 _3932_ (.A(_0627_),
    .B(_0633_),
    .C(_0638_),
    .D(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nand2_1 _3933_ (.A(_0421_),
    .B(_3030_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _3934_ (.A(_0425_),
    .B(_2932_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _3935_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__a221oi_1 _3936_ (.A1(_0415_),
    .A2(_3067_),
    .B1(_0418_),
    .B2(_0323_),
    .C1(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__buf_4 _3937_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .X(_0647_));
 sky130_fd_sc_hd__buf_4 _3938_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_0648_));
 sky130_fd_sc_hd__buf_4 _3939_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0649_));
 sky130_fd_sc_hd__nand2_1 _3940_ (.A(_0438_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__clkbuf_8 _3941_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _3942_ (.A(_0442_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _3943_ (.A(_0650_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__a221oi_1 _3944_ (.A1(_0647_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_0648_),
    .C1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__inv_2 _3945_ (.A(_2987_),
    .Y(_0655_));
 sky130_fd_sc_hd__inv_2 _3946_ (.A(_2839_),
    .Y(_0656_));
 sky130_fd_sc_hd__o22ai_1 _3947_ (.A1(_0655_),
    .A2(_0450_),
    .B1(_0656_),
    .B2(_0454_),
    .Y(_0657_));
 sky130_fd_sc_hd__a22o_1 _3948_ (.A1(_0456_),
    .A2(_0459_),
    .B1(_0458_),
    .B2(_2977_),
    .X(_0658_));
 sky130_fd_sc_hd__nor2_1 _3949_ (.A(_0657_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__inv_2 _3950_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _3951_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_0661_));
 sky130_fd_sc_hd__o22ai_1 _3952_ (.A1(_0660_),
    .A2(_0464_),
    .B1(_0661_),
    .B2(_0467_),
    .Y(_0662_));
 sky130_fd_sc_hd__a22o_1 _3953_ (.A1(_0469_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .B1(_0470_),
    .B2(_0439_),
    .X(_0663_));
 sky130_fd_sc_hd__nor2_1 _3954_ (.A(_0662_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__and4_1 _3955_ (.A(_0646_),
    .B(_0654_),
    .C(_0659_),
    .D(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__o22ai_1 _3956_ (.A1(_0492_),
    .A2(_0483_),
    .B1(_0346_),
    .B2(_0487_),
    .Y(_0666_));
 sky130_fd_sc_hd__a221oi_2 _3957_ (.A1(_0385_),
    .A2(_0478_),
    .B1(_0475_),
    .B2(_0480_),
    .C1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__o22ai_1 _3958_ (.A1(_0481_),
    .A2(_0491_),
    .B1(_0485_),
    .B2(_0493_),
    .Y(_0668_));
 sky130_fd_sc_hd__a22o_1 _3959_ (.A1(_0495_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .B1(_0496_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_0669_));
 sky130_fd_sc_hd__nor2_1 _3960_ (.A(_0668_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__inv_2 _3961_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_0671_));
 sky130_fd_sc_hd__o22ai_1 _3962_ (.A1(_0462_),
    .A2(_0500_),
    .B1(_0671_),
    .B2(_0503_),
    .Y(_0672_));
 sky130_fd_sc_hd__a22o_1 _3963_ (.A1(_0505_),
    .A2(_2786_),
    .B1(_0506_),
    .B2(_2777_),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_1 _3964_ (.A(_0672_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__inv_2 _3965_ (.A(_3053_),
    .Y(_0675_));
 sky130_fd_sc_hd__inv_2 _3966_ (.A(_3114_),
    .Y(_0676_));
 sky130_fd_sc_hd__o22ai_1 _3967_ (.A1(_0675_),
    .A2(_0512_),
    .B1(_0676_),
    .B2(_0515_),
    .Y(_0677_));
 sky130_fd_sc_hd__a22o_1 _3968_ (.A1(_0517_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .B1(_0518_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0678_));
 sky130_fd_sc_hd__nor2_1 _3969_ (.A(_0677_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__and4_1 _3970_ (.A(_0667_),
    .B(_0670_),
    .C(_0674_),
    .D(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__and4_1 _3971_ (.A(_0621_),
    .B(_0642_),
    .C(_0665_),
    .D(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__nand3_2 _3972_ (.A(_0602_),
    .B(_3113_),
    .C(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__o21a_1 _3973_ (.A1(_3078_),
    .A2(_0525_),
    .B1(_2776_),
    .X(_0683_));
 sky130_fd_sc_hd__a22o_1 _3974_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B1(_0682_),
    .B2(_0683_),
    .X(_0296_));
 sky130_fd_sc_hd__inv_2 _3975_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _3976_ (.A(_2837_),
    .B(_2904_),
    .Y(_0685_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(_2844_),
    .B(_2966_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _3978_ (.A(_0685_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__a221oi_2 _3979_ (.A1(_2921_),
    .A2(_2826_),
    .B1(_2886_),
    .B2(_2831_),
    .C1(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__a22o_1 _3980_ (.A1(_2853_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .B1(_2856_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_0689_));
 sky130_fd_sc_hd__a22o_1 _3981_ (.A1(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .A2(_2862_),
    .B1(_2864_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_0690_));
 sky130_fd_sc_hd__nor2_1 _3982_ (.A(_0689_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__inv_2 _3983_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _3984_ (.A(_2878_),
    .B(_2777_),
    .Y(_0693_));
 sky130_fd_sc_hd__o221a_1 _3985_ (.A1(_0671_),
    .A2(_2869_),
    .B1(_0692_),
    .B2(_2875_),
    .C1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_8 _3986_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(_2889_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__nand2_1 _3988_ (.A(_2893_),
    .B(_2804_),
    .Y(_0697_));
 sky130_fd_sc_hd__nand2_1 _3989_ (.A(_0696_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a221oi_1 _3990_ (.A1(_2884_),
    .A2(_2891_),
    .B1(_2887_),
    .B2(_2796_),
    .C1(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__and4_1 _3991_ (.A(_0688_),
    .B(_0691_),
    .C(_0694_),
    .D(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__o22ai_1 _3992_ (.A1(_2913_),
    .A2(_2910_),
    .B1(_0656_),
    .B2(_2915_),
    .Y(_0701_));
 sky130_fd_sc_hd__a221oi_1 _3993_ (.A1(_0447_),
    .A2(_2902_),
    .B1(_2987_),
    .B2(_2906_),
    .C1(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_1 _3994_ (.A(_2924_),
    .B(_2800_),
    .Y(_0703_));
 sky130_fd_sc_hd__nand2_1 _3995_ (.A(_2927_),
    .B(_2794_),
    .Y(_0704_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_0703_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__a221oi_1 _3997_ (.A1(_2919_),
    .A2(_2846_),
    .B1(_2922_),
    .B2(_2802_),
    .C1(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__buf_6 _3998_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_1 _3999_ (.A(_2943_),
    .B(_2792_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _4000_ (.A(_2947_),
    .B(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _4001_ (.A(_0708_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__a221oi_1 _4002_ (.A1(_0707_),
    .A2(_2938_),
    .B1(_2940_),
    .B2(_2798_),
    .C1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _4003_ (.A(_2960_),
    .B(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_0712_));
 sky130_fd_sc_hd__nand2_1 _4004_ (.A(_2964_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _4005_ (.A(_0712_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__a221oi_1 _4006_ (.A1(_0451_),
    .A2(_2954_),
    .B1(_0326_),
    .B2(_2958_),
    .C1(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__and4_1 _4007_ (.A(_0702_),
    .B(_0706_),
    .C(_0711_),
    .D(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__nand2_1 _4008_ (.A(_2985_),
    .B(_3009_),
    .Y(_0717_));
 sky130_fd_sc_hd__o21ai_1 _4009_ (.A1(_2991_),
    .A2(_2983_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a221oi_1 _4010_ (.A1(_0457_),
    .A2(_2975_),
    .B1(_2952_),
    .B2(_2980_),
    .C1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__or2_1 _4011_ (.A(_2982_),
    .B(_2994_),
    .X(_0720_));
 sky130_fd_sc_hd__nand2_1 _4012_ (.A(_2996_),
    .B(_0430_),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_1 _4013_ (.A(_3000_),
    .B(_0443_),
    .Y(_0722_));
 sky130_fd_sc_hd__o2111a_1 _4014_ (.A1(_3139_),
    .A2(_2992_),
    .B1(_0720_),
    .C1(_0721_),
    .D1(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__inv_2 _4015_ (.A(_3147_),
    .Y(_0724_));
 sky130_fd_sc_hd__inv_2 _4016_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_0725_));
 sky130_fd_sc_hd__o22ai_1 _4017_ (.A1(_0724_),
    .A2(_3015_),
    .B1(_0725_),
    .B2(_3021_),
    .Y(_0726_));
 sky130_fd_sc_hd__a221oi_1 _4018_ (.A1(_3013_),
    .A2(_3007_),
    .B1(_2956_),
    .B2(_3011_),
    .C1(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(_3034_),
    .B(_0651_),
    .Y(_0728_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_3038_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_0729_));
 sky130_fd_sc_hd__nand2_1 _4021_ (.A(_0728_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__a221oi_1 _4022_ (.A1(_3027_),
    .A2(_3030_),
    .B1(_3064_),
    .B2(_3032_),
    .C1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__and4_1 _4023_ (.A(_0719_),
    .B(_0723_),
    .C(_0727_),
    .D(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _4024_ (.A(_3051_),
    .B(_3058_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _4025_ (.A(_3056_),
    .B(_3114_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _4026_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__a221oi_2 _4027_ (.A1(_0513_),
    .A2(_3046_),
    .B1(_3048_),
    .B2(_0623_),
    .C1(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _4028_ (.A(_3068_),
    .B(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(_3071_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _4030_ (.A(_0737_),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__a221oi_1 _4031_ (.A1(_3062_),
    .A2(_2932_),
    .B1(_3065_),
    .B2(_0419_),
    .C1(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__inv_2 _4032_ (.A(_0459_),
    .Y(_0741_));
 sky130_fd_sc_hd__nand2_1 _4033_ (.A(_3087_),
    .B(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0742_));
 sky130_fd_sc_hd__o21ai_1 _4034_ (.A1(_0741_),
    .A2(_3085_),
    .B1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__a221oi_1 _4035_ (.A1(_3076_),
    .A2(_0591_),
    .B1(_0479_),
    .B2(_3081_),
    .C1(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__clkbuf_8 _4036_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_8 _4037_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_0746_));
 sky130_fd_sc_hd__nand2_1 _4038_ (.A(_3099_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _4039_ (.A(_3102_),
    .B(_0631_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _4040_ (.A(_0747_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__a221oi_1 _4041_ (.A1(_0745_),
    .A2(_3094_),
    .B1(_3096_),
    .B2(_0746_),
    .C1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__and4_1 _4042_ (.A(_0736_),
    .B(_0740_),
    .C(_0744_),
    .D(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__and4_1 _4043_ (.A(_0700_),
    .B(_0716_),
    .C(_0732_),
    .D(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__nand2_1 _4044_ (.A(_3125_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0753_));
 sky130_fd_sc_hd__o21ai_1 _4045_ (.A1(_0618_),
    .A2(_3123_),
    .B1(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__a221oi_1 _4046_ (.A1(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .A2(_3116_),
    .B1(_0391_),
    .B2(_3120_),
    .C1(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__or2_1 _4047_ (.A(_3084_),
    .B(_3136_),
    .X(_0756_));
 sky130_fd_sc_hd__or2_1 _4048_ (.A(_3135_),
    .B(_3140_),
    .X(_0757_));
 sky130_fd_sc_hd__nand2_1 _4049_ (.A(_3143_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0758_));
 sky130_fd_sc_hd__o2111a_1 _4050_ (.A1(_3122_),
    .A2(_3132_),
    .B1(_0756_),
    .C1(_0757_),
    .D1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nand2_1 _4051_ (.A(_0324_),
    .B(_0338_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _4052_ (.A(_0328_),
    .B(_2971_),
    .Y(_0761_));
 sky130_fd_sc_hd__nand2_1 _4053_ (.A(_0760_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__a221oi_2 _4054_ (.A1(_3017_),
    .A2(_3149_),
    .B1(_3151_),
    .B2(_0352_),
    .C1(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__inv_2 _4055_ (.A(_3118_),
    .Y(_0764_));
 sky130_fd_sc_hd__o22ai_1 _4056_ (.A1(_0764_),
    .A2(_0343_),
    .B1(_0675_),
    .B2(_0347_),
    .Y(_0765_));
 sky130_fd_sc_hd__a221oi_1 _4057_ (.A1(_3050_),
    .A2(_0336_),
    .B1(_0384_),
    .B2(_0340_),
    .C1(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__and4_1 _4058_ (.A(_0755_),
    .B(_0759_),
    .C(_0763_),
    .D(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_8 _4059_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_0768_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(_0359_),
    .B(_0364_),
    .Y(_0769_));
 sky130_fd_sc_hd__nand2_1 _4061_ (.A(_0362_),
    .B(_3079_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _4062_ (.A(_0769_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__a221oi_1 _4063_ (.A1(_3029_),
    .A2(_0354_),
    .B1(_0356_),
    .B2(_0768_),
    .C1(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__or2b_1 _4064_ (.A(_0368_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0773_));
 sky130_fd_sc_hd__nand2_1 _4065_ (.A(_0371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0774_));
 sky130_fd_sc_hd__nand2_1 _4066_ (.A(_0374_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_1 _4067_ (.A(_0377_),
    .B(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_0776_));
 sky130_fd_sc_hd__and4_1 _4068_ (.A(_0773_),
    .B(_0774_),
    .C(_0775_),
    .D(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _4069_ (.A(_0389_),
    .B(_0395_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand2_1 _4070_ (.A(_0393_),
    .B(_0475_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _4071_ (.A(_0778_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__a221oi_1 _4072_ (.A1(_0382_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .B1(_0416_),
    .B2(_0387_),
    .C1(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__a22o_1 _4073_ (.A1(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .A2(_0400_),
    .B1(_0403_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_1 _4074_ (.A1(_0406_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .B1(_0408_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0783_));
 sky130_fd_sc_hd__nor2_1 _4075_ (.A(_0782_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__and4_1 _4076_ (.A(_0772_),
    .B(_0777_),
    .C(_0781_),
    .D(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _4077_ (.A(_0421_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _4078_ (.A(_0425_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0787_));
 sky130_fd_sc_hd__nand2_1 _4079_ (.A(_0786_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__a221oi_1 _4080_ (.A1(_0415_),
    .A2(_0584_),
    .B1(_0418_),
    .B2(_0613_),
    .C1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2_1 _4081_ (.A(_0437_),
    .B(_3002_),
    .Y(_0790_));
 sky130_fd_sc_hd__buf_4 _4082_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .X(_0791_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(_0441_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_1 _4084_ (.A(_0790_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__a221oi_1 _4085_ (.A1(_0330_),
    .A2(_0432_),
    .B1(_0434_),
    .B2(_2998_),
    .C1(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _4086_ (.A(_3005_),
    .Y(_0795_));
 sky130_fd_sc_hd__inv_2 _4087_ (.A(_2899_),
    .Y(_0796_));
 sky130_fd_sc_hd__o22ai_1 _4088_ (.A1(_0795_),
    .A2(_0449_),
    .B1(_0796_),
    .B2(_0453_),
    .Y(_0797_));
 sky130_fd_sc_hd__a22o_1 _4089_ (.A1(_0456_),
    .A2(_2977_),
    .B1(_0458_),
    .B2(_2908_),
    .X(_0798_));
 sky130_fd_sc_hd__nor2_1 _4090_ (.A(_0797_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__inv_2 _4091_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_0800_));
 sky130_fd_sc_hd__inv_2 _4092_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_0801_));
 sky130_fd_sc_hd__o22ai_1 _4093_ (.A1(_0800_),
    .A2(_0463_),
    .B1(_0801_),
    .B2(_0466_),
    .Y(_0802_));
 sky130_fd_sc_hd__a22o_1 _4094_ (.A1(_0469_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .B1(_0470_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0803_));
 sky130_fd_sc_hd__nor2_1 _4095_ (.A(_0802_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__and4_1 _4096_ (.A(_0789_),
    .B(_0794_),
    .C(_0799_),
    .D(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__o22ai_1 _4097_ (.A1(_0485_),
    .A2(_0482_),
    .B1(_0511_),
    .B2(_0486_),
    .Y(_0806_));
 sky130_fd_sc_hd__a221oi_1 _4098_ (.A1(_0634_),
    .A2(_0477_),
    .B1(_0385_),
    .B2(_2757_),
    .C1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__o22ai_1 _4099_ (.A1(_0492_),
    .A2(_0491_),
    .B1(_0346_),
    .B2(_0493_),
    .Y(_0808_));
 sky130_fd_sc_hd__a22o_1 _4100_ (.A1(_0495_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .B1(_0496_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0809_));
 sky130_fd_sc_hd__nor2_1 _4101_ (.A(_0808_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_2 _4102_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_0811_));
 sky130_fd_sc_hd__o22ai_1 _4103_ (.A1(_0660_),
    .A2(_0500_),
    .B1(_0811_),
    .B2(_0502_),
    .Y(_0812_));
 sky130_fd_sc_hd__a22o_1 _4104_ (.A1(_0505_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .B1(_0506_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_1 _4105_ (.A(_0812_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _4106_ (.A(_3044_),
    .Y(_0815_));
 sky130_fd_sc_hd__inv_2 _4107_ (.A(_3127_),
    .Y(_0816_));
 sky130_fd_sc_hd__o22ai_1 _4108_ (.A1(_0815_),
    .A2(_0512_),
    .B1(_0816_),
    .B2(_0515_),
    .Y(_0817_));
 sky130_fd_sc_hd__a22o_1 _4109_ (.A1(_0517_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .B1(_0518_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0818_));
 sky130_fd_sc_hd__nor2_1 _4110_ (.A(_0817_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__and4_1 _4111_ (.A(_0807_),
    .B(_0810_),
    .C(_0814_),
    .D(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__and4_1 _4112_ (.A(_0767_),
    .B(_0785_),
    .C(_0805_),
    .D(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__o21ai_1 _4113_ (.A1(_0589_),
    .A2(_3112_),
    .B1(_2775_),
    .Y(_0822_));
 sky130_fd_sc_hd__a31o_1 _4114_ (.A1(_0752_),
    .A2(_0821_),
    .A3(_0525_),
    .B1(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__o21ai_1 _4115_ (.A1(_2776_),
    .A2(_0684_),
    .B1(_0823_),
    .Y(_0295_));
 sky130_fd_sc_hd__clkbuf_4 _4116_ (.A(_2862_),
    .X(_0824_));
 sky130_fd_sc_hd__clkbuf_4 _4117_ (.A(_2864_),
    .X(_0825_));
 sky130_fd_sc_hd__a22o_1 _4118_ (.A1(_2854_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .B1(_2857_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_0826_));
 sky130_fd_sc_hd__a221oi_1 _4119_ (.A1(_0524_),
    .A2(_0824_),
    .B1(_2846_),
    .B2(_0825_),
    .C1(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__nand2_1 _4120_ (.A(_2838_),
    .B(_0447_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _4121_ (.A(_2845_),
    .B(_2891_),
    .Y(_0829_));
 sky130_fd_sc_hd__nand2_1 _4122_ (.A(_0828_),
    .B(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__a221oi_2 _4123_ (.A1(_2828_),
    .A2(_2827_),
    .B1(_2966_),
    .B2(_2832_),
    .C1(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__inv_2 _4124_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_1 _4125_ (.A(_2879_),
    .B(_2786_),
    .Y(_0833_));
 sky130_fd_sc_hd__o221a_1 _4126_ (.A1(_0811_),
    .A2(_2870_),
    .B1(_0832_),
    .B2(_2875_),
    .C1(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__nand2_1 _4127_ (.A(_2890_),
    .B(_2880_),
    .Y(_0835_));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(_2894_),
    .B(_2806_),
    .Y(_0836_));
 sky130_fd_sc_hd__nand2_1 _4129_ (.A(_0835_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__a221oi_1 _4130_ (.A1(_2885_),
    .A2(_0537_),
    .B1(_2888_),
    .B2(_2798_),
    .C1(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__and4_1 _4131_ (.A(_0827_),
    .B(_0831_),
    .C(_0834_),
    .D(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o22ai_1 _4132_ (.A1(_0452_),
    .A2(_2911_),
    .B1(_0796_),
    .B2(_2916_),
    .Y(_0840_));
 sky130_fd_sc_hd__a221oi_1 _4133_ (.A1(_2987_),
    .A2(_2903_),
    .B1(_3005_),
    .B2(_2907_),
    .C1(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__nand2_1 _4134_ (.A(_2925_),
    .B(_2802_),
    .Y(_0842_));
 sky130_fd_sc_hd__nand2_1 _4135_ (.A(_2928_),
    .B(_2796_),
    .Y(_0843_));
 sky130_fd_sc_hd__nand2_1 _4136_ (.A(_0842_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__a221oi_2 _4137_ (.A1(_2920_),
    .A2(_2886_),
    .B1(_2923_),
    .B2(_2804_),
    .C1(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _4138_ (.A(_2944_),
    .B(_2794_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _4139_ (.A(_2948_),
    .B(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _4140_ (.A(_0846_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__a221oi_1 _4141_ (.A1(_3098_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2800_),
    .C1(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_1 _4142_ (.A(_2961_),
    .B(_2921_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _4143_ (.A(_2965_),
    .B(_0695_),
    .Y(_0851_));
 sky130_fd_sc_hd__nand2_1 _4144_ (.A(_0850_),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__a221oi_1 _4145_ (.A1(_2839_),
    .A2(_2955_),
    .B1(_3017_),
    .B2(_2959_),
    .C1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__and4_1 _4146_ (.A(_0841_),
    .B(_0845_),
    .C(_0849_),
    .D(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _4147_ (.A(_2986_),
    .B(_3013_),
    .Y(_0855_));
 sky130_fd_sc_hd__o21ai_1 _4148_ (.A1(_0564_),
    .A2(_2984_),
    .B1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a221oi_1 _4149_ (.A1(_0459_),
    .A2(_2976_),
    .B1(_2912_),
    .B2(_2981_),
    .C1(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__buf_2 _4150_ (.A(_2994_),
    .X(_0858_));
 sky130_fd_sc_hd__or2_1 _4151_ (.A(_0560_),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__nand2_1 _4152_ (.A(_2997_),
    .B(_0647_),
    .Y(_0860_));
 sky130_fd_sc_hd__nand2_1 _4153_ (.A(_3001_),
    .B(_0651_),
    .Y(_0861_));
 sky130_fd_sc_hd__o2111a_1 _4154_ (.A1(_0609_),
    .A2(_2993_),
    .B1(_0859_),
    .C1(_0860_),
    .D1(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__inv_2 _4155_ (.A(_0326_),
    .Y(_0863_));
 sky130_fd_sc_hd__inv_2 _4156_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_0864_));
 sky130_fd_sc_hd__o22ai_1 _4157_ (.A1(_0863_),
    .A2(_3016_),
    .B1(_0864_),
    .B2(_3022_),
    .Y(_0865_));
 sky130_fd_sc_hd__a221oi_1 _4158_ (.A1(_2956_),
    .A2(_3008_),
    .B1(_3147_),
    .B2(_3012_),
    .C1(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(_3035_),
    .B(_0791_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand2_1 _4160_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_0868_));
 sky130_fd_sc_hd__nand2_1 _4161_ (.A(_0867_),
    .B(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__a221oi_1 _4162_ (.A1(_3028_),
    .A2(_0574_),
    .B1(_0426_),
    .B2(_3033_),
    .C1(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__and4_1 _4163_ (.A(_0857_),
    .B(_0862_),
    .C(_0866_),
    .D(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__nand2_1 _4164_ (.A(_3052_),
    .B(_0513_),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_1 _4165_ (.A(_3057_),
    .B(_3127_),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _4166_ (.A(_0872_),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__a221oi_1 _4167_ (.A1(_3114_),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0768_),
    .C1(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _4168_ (.A(_3069_),
    .B(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_0876_));
 sky130_fd_sc_hd__nand2_1 _4169_ (.A(_3072_),
    .B(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_0877_));
 sky130_fd_sc_hd__nand2_1 _4170_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__a221oi_1 _4171_ (.A1(_3063_),
    .A2(_0550_),
    .B1(_3066_),
    .B2(_0323_),
    .C1(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__inv_2 _4172_ (.A(_2977_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _4173_ (.A(_3088_),
    .B(_0648_),
    .Y(_0881_));
 sky130_fd_sc_hd__o21ai_1 _4174_ (.A1(_0880_),
    .A2(_3086_),
    .B1(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__a221oi_1 _4175_ (.A1(_3077_),
    .A2(_0436_),
    .B1(_0475_),
    .B2(_3082_),
    .C1(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__clkbuf_8 _4176_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_0884_));
 sky130_fd_sc_hd__nand2_1 _4177_ (.A(_3100_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_0885_));
 sky130_fd_sc_hd__nand2_1 _4178_ (.A(_3103_),
    .B(_0471_),
    .Y(_0886_));
 sky130_fd_sc_hd__nand2_1 _4179_ (.A(_0885_),
    .B(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__a221oi_1 _4180_ (.A1(_0884_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0410_),
    .C1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__and4_2 _4181_ (.A(_0875_),
    .B(_0879_),
    .C(_0883_),
    .D(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__and4_1 _4182_ (.A(_0839_),
    .B(_0854_),
    .C(_0871_),
    .D(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__nand2_1 _4183_ (.A(_3126_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_0891_));
 sky130_fd_sc_hd__o21ai_1 _4184_ (.A1(_0764_),
    .A2(_3124_),
    .B1(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__a221oi_2 _4185_ (.A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .A2(_3117_),
    .B1(_3079_),
    .B2(_3121_),
    .C1(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__or2_1 _4186_ (.A(_0590_),
    .B(_3137_),
    .X(_0894_));
 sky130_fd_sc_hd__or2_1 _4187_ (.A(_0607_),
    .B(_3141_),
    .X(_0895_));
 sky130_fd_sc_hd__nand2_1 _4188_ (.A(_3144_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0896_));
 sky130_fd_sc_hd__o2111a_1 _4189_ (.A1(_0342_),
    .A2(_3133_),
    .B1(_0894_),
    .C1(_0895_),
    .D1(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _4190_ (.A(_0325_),
    .B(_0334_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_1 _4191_ (.A(_0329_),
    .B(_3083_),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _4192_ (.A(_0898_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__a221oi_1 _4193_ (.A1(_0338_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0622_),
    .C1(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__inv_2 _4194_ (.A(_0364_),
    .Y(_0902_));
 sky130_fd_sc_hd__o22ai_1 _4195_ (.A1(_0902_),
    .A2(_0344_),
    .B1(_0815_),
    .B2(_0348_),
    .Y(_0903_));
 sky130_fd_sc_hd__a221oi_1 _4196_ (.A1(_0358_),
    .A2(_0337_),
    .B1(_3050_),
    .B2(_0341_),
    .C1(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__and4_1 _4197_ (.A(_0893_),
    .B(_0897_),
    .C(_0901_),
    .D(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_4 _4198_ (.A(_0495_),
    .X(_0906_));
 sky130_fd_sc_hd__clkbuf_4 _4199_ (.A(_0496_),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_4 _4200_ (.A(_0491_),
    .X(_0908_));
 sky130_fd_sc_hd__clkbuf_4 _4201_ (.A(_0493_),
    .X(_0909_));
 sky130_fd_sc_hd__o22ai_1 _4202_ (.A1(_0485_),
    .A2(_0908_),
    .B1(_0511_),
    .B2(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__a221oi_1 _4203_ (.A1(_0595_),
    .A2(_0906_),
    .B1(_0745_),
    .B2(_0907_),
    .C1(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__o22ai_1 _4204_ (.A1(_0346_),
    .A2(_0483_),
    .B1(_0675_),
    .B2(_0487_),
    .Y(_0912_));
 sky130_fd_sc_hd__a221oi_1 _4205_ (.A1(_0416_),
    .A2(_0478_),
    .B1(_0634_),
    .B2(_0480_),
    .C1(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__inv_2 _4206_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_0914_));
 sky130_fd_sc_hd__clkbuf_4 _4207_ (.A(_0500_),
    .X(_0915_));
 sky130_fd_sc_hd__o22ai_1 _4208_ (.A1(_0914_),
    .A2(_0503_),
    .B1(_0800_),
    .B2(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__buf_4 _4209_ (.A(_0505_),
    .X(_0917_));
 sky130_fd_sc_hd__buf_4 _4210_ (.A(_0506_),
    .X(_0918_));
 sky130_fd_sc_hd__a22o_1 _4211_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .B1(_0918_),
    .B2(_2788_),
    .X(_0919_));
 sky130_fd_sc_hd__nor2_1 _4212_ (.A(_0916_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__inv_2 _4213_ (.A(_3058_),
    .Y(_0921_));
 sky130_fd_sc_hd__clkbuf_4 _4214_ (.A(_0512_),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_4 _4215_ (.A(_0515_),
    .X(_0923_));
 sky130_fd_sc_hd__o22ai_1 _4216_ (.A1(_0921_),
    .A2(_0922_),
    .B1(_3131_),
    .B2(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__clkbuf_4 _4217_ (.A(_0517_),
    .X(_0925_));
 sky130_fd_sc_hd__clkbuf_4 _4218_ (.A(_0518_),
    .X(_0926_));
 sky130_fd_sc_hd__a22o_1 _4219_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .B1(_0926_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_0927_));
 sky130_fd_sc_hd__nor2_1 _4220_ (.A(_0924_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__and4_1 _4221_ (.A(_0911_),
    .B(_0913_),
    .C(_0920_),
    .D(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_4 _4222_ (.A(_0456_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_4 _4223_ (.A(_0458_),
    .X(_0931_));
 sky130_fd_sc_hd__inv_2 _4224_ (.A(_3009_),
    .Y(_0932_));
 sky130_fd_sc_hd__inv_2 _4225_ (.A(_2904_),
    .Y(_0933_));
 sky130_fd_sc_hd__o22ai_1 _4226_ (.A1(_0932_),
    .A2(_0450_),
    .B1(_0933_),
    .B2(_0454_),
    .Y(_0934_));
 sky130_fd_sc_hd__a221oi_1 _4227_ (.A1(_2908_),
    .A2(_0930_),
    .B1(_2952_),
    .B2(_0931_),
    .C1(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__clkbuf_4 _4228_ (.A(_0469_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_4 _4229_ (.A(_0470_),
    .X(_0937_));
 sky130_fd_sc_hd__inv_2 _4230_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_0938_));
 sky130_fd_sc_hd__inv_2 _4231_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_0939_));
 sky130_fd_sc_hd__o22ai_1 _4232_ (.A1(_0938_),
    .A2(_0464_),
    .B1(_0939_),
    .B2(_0467_),
    .Y(_0940_));
 sky130_fd_sc_hd__a221oi_1 _4233_ (.A1(_0649_),
    .A2(_0936_),
    .B1(_3002_),
    .B2(_0937_),
    .C1(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__nand2_1 _4234_ (.A(_0438_),
    .B(_3036_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _4235_ (.A(_0442_),
    .B(_2962_),
    .Y(_0943_));
 sky130_fd_sc_hd__nand2_1 _4236_ (.A(_0942_),
    .B(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__a221oi_1 _4237_ (.A1(_3134_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_0566_),
    .C1(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__nand2_1 _4238_ (.A(_0421_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_1 _4239_ (.A(_0425_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _4240_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__a221oi_1 _4241_ (.A1(_0415_),
    .A2(_0419_),
    .B1(_0418_),
    .B2(_0352_),
    .C1(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__and4_1 _4242_ (.A(_0935_),
    .B(_0941_),
    .C(_0945_),
    .D(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(_0360_),
    .B(_0391_),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _4244_ (.A(_0363_),
    .B(_0395_),
    .Y(_0952_));
 sky130_fd_sc_hd__nand2_1 _4245_ (.A(_0951_),
    .B(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__a221oi_1 _4246_ (.A1(_0422_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_3092_),
    .C1(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__nand2b_1 _4247_ (.A_N(_0369_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _4248_ (.A(_0372_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0956_));
 sky130_fd_sc_hd__nand2_1 _4249_ (.A(_0375_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0957_));
 sky130_fd_sc_hd__nand2_1 _4250_ (.A(_0378_),
    .B(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_0958_));
 sky130_fd_sc_hd__and4_1 _4251_ (.A(_0955_),
    .B(_0956_),
    .C(_0957_),
    .D(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__nand2_1 _4252_ (.A(_0390_),
    .B(_0479_),
    .Y(_0960_));
 sky130_fd_sc_hd__nand2_1 _4253_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_0961_));
 sky130_fd_sc_hd__nand2_1 _4254_ (.A(_0960_),
    .B(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__a221oi_1 _4255_ (.A1(_0383_),
    .A2(_0623_),
    .B1(_3067_),
    .B2(_0388_),
    .C1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__a22o_1 _4256_ (.A1(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_0964_));
 sky130_fd_sc_hd__a22o_1 _4257_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .B1(_0409_),
    .B2(_0631_),
    .X(_0965_));
 sky130_fd_sc_hd__nor2_1 _4258_ (.A(_0964_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__and4_1 _4259_ (.A(_0954_),
    .B(_0959_),
    .C(_0963_),
    .D(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__and4_1 _4260_ (.A(_0905_),
    .B(_0929_),
    .C(_0950_),
    .D(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__nand3_2 _4261_ (.A(_0890_),
    .B(_3113_),
    .C(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__o21a_1 _4262_ (.A1(_0591_),
    .A2(_0525_),
    .B1(_2776_),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _4263_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B1(_0969_),
    .B2(_0970_),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_1 _4264_ (.A1(_2854_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .B1(_2857_),
    .B2(_2814_),
    .X(_0971_));
 sky130_fd_sc_hd__a221oi_1 _4265_ (.A1(_3078_),
    .A2(_0824_),
    .B1(_2886_),
    .B2(_0825_),
    .C1(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__nand2_1 _4266_ (.A(_2838_),
    .B(_2987_),
    .Y(_0973_));
 sky130_fd_sc_hd__nand2_1 _4267_ (.A(_2845_),
    .B(_0537_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_1 _4268_ (.A(_0973_),
    .B(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__a221oi_2 _4269_ (.A1(_2846_),
    .A2(_2827_),
    .B1(_2891_),
    .B2(_2832_),
    .C1(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__inv_2 _4270_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_0977_));
 sky130_fd_sc_hd__nand2_1 _4271_ (.A(_2879_),
    .B(_2788_),
    .Y(_0978_));
 sky130_fd_sc_hd__o221a_1 _4272_ (.A1(_0914_),
    .A2(_2870_),
    .B1(_0977_),
    .B2(_2875_),
    .C1(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__nand2_1 _4273_ (.A(_2890_),
    .B(_0507_),
    .Y(_0980_));
 sky130_fd_sc_hd__nand2_1 _4274_ (.A(_2894_),
    .B(_2808_),
    .Y(_0981_));
 sky130_fd_sc_hd__nand2_1 _4275_ (.A(_0980_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__a221oi_1 _4276_ (.A1(_2885_),
    .A2(_0695_),
    .B1(_2888_),
    .B2(_2800_),
    .C1(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__and4_1 _4277_ (.A(_0972_),
    .B(_0976_),
    .C(_0979_),
    .D(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__o22ai_1 _4278_ (.A1(_0656_),
    .A2(_2911_),
    .B1(_0933_),
    .B2(_2916_),
    .Y(_0985_));
 sky130_fd_sc_hd__a221oi_1 _4279_ (.A1(_3005_),
    .A2(_2903_),
    .B1(_3009_),
    .B2(_2907_),
    .C1(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__nand2_1 _4280_ (.A(_2925_),
    .B(_2804_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand2_1 _4281_ (.A(_2928_),
    .B(_2798_),
    .Y(_0988_));
 sky130_fd_sc_hd__nand2_1 _4282_ (.A(_0987_),
    .B(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__a221oi_1 _4283_ (.A1(_2920_),
    .A2(_2966_),
    .B1(_2923_),
    .B2(_2806_),
    .C1(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_2944_),
    .B(_2796_),
    .Y(_0991_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_2948_),
    .B(_2812_),
    .Y(_0992_));
 sky130_fd_sc_hd__nand2_1 _4286_ (.A(_0991_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__a221oi_1 _4287_ (.A1(_0596_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2802_),
    .C1(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand2_1 _4288_ (.A(_2961_),
    .B(_2828_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _4289_ (.A(_2965_),
    .B(_2880_),
    .Y(_0996_));
 sky130_fd_sc_hd__nand2_1 _4290_ (.A(_0995_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__a221oi_1 _4291_ (.A1(_2899_),
    .A2(_2955_),
    .B1(_0338_),
    .B2(_2959_),
    .C1(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__and4_1 _4292_ (.A(_0986_),
    .B(_0990_),
    .C(_0994_),
    .D(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(_2986_),
    .B(_2956_),
    .Y(_1000_));
 sky130_fd_sc_hd__o21ai_1 _4294_ (.A1(_3139_),
    .A2(_2984_),
    .B1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__a221oi_1 _4295_ (.A1(_2977_),
    .A2(_2976_),
    .B1(_0451_),
    .B2(_2981_),
    .C1(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__or2_1 _4296_ (.A(_2991_),
    .B(_0858_),
    .X(_1003_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(_2997_),
    .B(_0330_),
    .Y(_1004_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_3001_),
    .B(_0791_),
    .Y(_1005_));
 sky130_fd_sc_hd__o2111a_1 _4299_ (.A1(_3135_),
    .A2(_2993_),
    .B1(_1003_),
    .C1(_1004_),
    .D1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__inv_2 _4300_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_1007_));
 sky130_fd_sc_hd__o22ai_1 _4301_ (.A1(_3018_),
    .A2(_3016_),
    .B1(_1007_),
    .B2(_3022_),
    .Y(_1008_));
 sky130_fd_sc_hd__a221oi_1 _4302_ (.A1(_3147_),
    .A2(_3008_),
    .B1(_0326_),
    .B2(_3012_),
    .C1(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__nand2_1 _4303_ (.A(_3035_),
    .B(_2962_),
    .Y(_1010_));
 sky130_fd_sc_hd__nand2_1 _4304_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1011_));
 sky130_fd_sc_hd__nand2_1 _4305_ (.A(_1010_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__a221oi_1 _4306_ (.A1(_3028_),
    .A2(_3064_),
    .B1(_2932_),
    .B2(_3033_),
    .C1(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__and4_1 _4307_ (.A(_1002_),
    .B(_1006_),
    .C(_1009_),
    .D(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__nand2_1 _4308_ (.A(_3052_),
    .B(_3114_),
    .Y(_1015_));
 sky130_fd_sc_hd__nand2_1 _4309_ (.A(_3057_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1016_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(_1015_),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__a221oi_1 _4311_ (.A1(_3127_),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_3092_),
    .C1(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_3069_),
    .B(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .Y(_1019_));
 sky130_fd_sc_hd__nand2_1 _4313_ (.A(_3072_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_1020_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_1019_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__a221oi_1 _4315_ (.A1(_3063_),
    .A2(_0707_),
    .B1(_3066_),
    .B2(_0613_),
    .C1(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2_1 _4316_ (.A(_3088_),
    .B(_2998_),
    .Y(_1023_));
 sky130_fd_sc_hd__o21ai_1 _4317_ (.A1(_2909_),
    .A2(_3086_),
    .B1(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__a221oi_1 _4318_ (.A1(_3077_),
    .A2(_0648_),
    .B1(_0385_),
    .B2(_3082_),
    .C1(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand2_1 _4319_ (.A(_3100_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1026_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(_3103_),
    .B(_0439_),
    .Y(_1027_));
 sky130_fd_sc_hd__nand2_1 _4321_ (.A(_1026_),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__a221oi_1 _4322_ (.A1(_0484_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_3104_),
    .C1(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__and4_1 _4323_ (.A(_1018_),
    .B(_1022_),
    .C(_1025_),
    .D(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__and4_1 _4324_ (.A(_0984_),
    .B(_0999_),
    .C(_1014_),
    .D(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(_3126_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1032_));
 sky130_fd_sc_hd__o21ai_1 _4326_ (.A1(_0902_),
    .A2(_3124_),
    .B1(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__a221oi_1 _4327_ (.A1(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .A2(_3117_),
    .B1(_0395_),
    .B2(_3121_),
    .C1(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__or2_1 _4328_ (.A(_0741_),
    .B(_3137_),
    .X(_1035_));
 sky130_fd_sc_hd__or2_1 _4329_ (.A(_3084_),
    .B(_3141_),
    .X(_1036_));
 sky130_fd_sc_hd__nand2_1 _4330_ (.A(_3144_),
    .B(_3118_),
    .Y(_1037_));
 sky130_fd_sc_hd__o2111a_1 _4331_ (.A1(_0618_),
    .A2(_3133_),
    .B1(_1035_),
    .C1(_1036_),
    .D1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_0325_),
    .B(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(_0329_),
    .B(_0457_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_1039_),
    .B(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__a221oi_1 _4335_ (.A1(_0334_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_3029_),
    .C1(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__inv_2 _4336_ (.A(_0391_),
    .Y(_1043_));
 sky130_fd_sc_hd__o22ai_1 _4337_ (.A1(_1043_),
    .A2(_0344_),
    .B1(_0921_),
    .B2(_0348_),
    .Y(_1044_));
 sky130_fd_sc_hd__a221oi_1 _4338_ (.A1(_0623_),
    .A2(_0337_),
    .B1(_0358_),
    .B2(_0341_),
    .C1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__and4_1 _4339_ (.A(_1034_),
    .B(_1038_),
    .C(_1042_),
    .D(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__o22ai_1 _4340_ (.A1(_0346_),
    .A2(_0908_),
    .B1(_0675_),
    .B2(_0909_),
    .Y(_1047_));
 sky130_fd_sc_hd__a221oi_1 _4341_ (.A1(_0745_),
    .A2(_0906_),
    .B1(_0884_),
    .B2(_0907_),
    .C1(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__o22ai_1 _4342_ (.A1(_0511_),
    .A2(_0483_),
    .B1(_0815_),
    .B2(_0487_),
    .Y(_1049_));
 sky130_fd_sc_hd__a221oi_1 _4343_ (.A1(_3067_),
    .A2(_0478_),
    .B1(_0416_),
    .B2(_0480_),
    .C1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__o22ai_1 _4344_ (.A1(_2871_),
    .A2(_0503_),
    .B1(_0938_),
    .B2(_0915_),
    .Y(_1051_));
 sky130_fd_sc_hd__a22o_1 _4345_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .B1(_0918_),
    .B2(_2790_),
    .X(_1052_));
 sky130_fd_sc_hd__nor2_1 _4346_ (.A(_1051_),
    .B(_1052_),
    .Y(_1053_));
 sky130_fd_sc_hd__o22ai_1 _4347_ (.A1(_0514_),
    .A2(_0922_),
    .B1(_0606_),
    .B2(_0923_),
    .Y(_1054_));
 sky130_fd_sc_hd__a22o_1 _4348_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .B1(_0926_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_1055_));
 sky130_fd_sc_hd__nor2_1 _4349_ (.A(_1054_),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__and4_1 _4350_ (.A(_1048_),
    .B(_1050_),
    .C(_1053_),
    .D(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__o22ai_1 _4351_ (.A1(_3014_),
    .A2(_0450_),
    .B1(_0448_),
    .B2(_0454_),
    .Y(_1058_));
 sky130_fd_sc_hd__a221oi_1 _4352_ (.A1(_2952_),
    .A2(_0930_),
    .B1(_2912_),
    .B2(_0931_),
    .C1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__inv_2 _4353_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_1060_));
 sky130_fd_sc_hd__o22ai_1 _4354_ (.A1(_1060_),
    .A2(_0464_),
    .B1(_0499_),
    .B2(_0467_),
    .Y(_1061_));
 sky130_fd_sc_hd__a221oi_1 _4355_ (.A1(_3002_),
    .A2(_0936_),
    .B1(_3036_),
    .B2(_0937_),
    .C1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_0438_),
    .B(_0443_),
    .Y(_1063_));
 sky130_fd_sc_hd__nand2_1 _4357_ (.A(_0442_),
    .B(_2817_),
    .Y(_1064_));
 sky130_fd_sc_hd__nand2_1 _4358_ (.A(_1063_),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__a221oi_1 _4359_ (.A1(_2971_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_0430_),
    .C1(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(_0421_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1067_));
 sky130_fd_sc_hd__nand2_1 _4361_ (.A(_0425_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_1068_));
 sky130_fd_sc_hd__nand2_1 _4362_ (.A(_1067_),
    .B(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__a221oi_1 _4363_ (.A1(_0415_),
    .A2(_0323_),
    .B1(_0418_),
    .B2(_0622_),
    .C1(_1069_),
    .Y(_1070_));
 sky130_fd_sc_hd__and4_1 _4364_ (.A(_1059_),
    .B(_1062_),
    .C(_1066_),
    .D(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(_0360_),
    .B(_3079_),
    .Y(_1072_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(_0363_),
    .B(_0479_),
    .Y(_1073_));
 sky130_fd_sc_hd__nand2_1 _4367_ (.A(_1072_),
    .B(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__a221oi_2 _4368_ (.A1(_3030_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0595_),
    .C1(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__nand2b_1 _4369_ (.A_N(_0369_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_1076_));
 sky130_fd_sc_hd__nand2_1 _4370_ (.A(_0372_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_1077_));
 sky130_fd_sc_hd__nand2_1 _4371_ (.A(_0375_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1078_));
 sky130_fd_sc_hd__nand2_1 _4372_ (.A(_0378_),
    .B(_0649_),
    .Y(_1079_));
 sky130_fd_sc_hd__and4_1 _4373_ (.A(_1076_),
    .B(_1077_),
    .C(_1078_),
    .D(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__nand2_1 _4374_ (.A(_0390_),
    .B(_0475_),
    .Y(_1081_));
 sky130_fd_sc_hd__nand2_1 _4375_ (.A(_0394_),
    .B(_0634_),
    .Y(_1082_));
 sky130_fd_sc_hd__nand2_1 _4376_ (.A(_1081_),
    .B(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__a221oi_1 _4377_ (.A1(_0383_),
    .A2(_0768_),
    .B1(_0584_),
    .B2(_0388_),
    .C1(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__a22o_1 _4378_ (.A1(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_1085_));
 sky130_fd_sc_hd__a22o_1 _4379_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .B1(_0409_),
    .B2(_0471_),
    .X(_1086_));
 sky130_fd_sc_hd__nor2_1 _4380_ (.A(_1085_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__and4_1 _4381_ (.A(_1075_),
    .B(_1080_),
    .C(_1084_),
    .D(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__and4_1 _4382_ (.A(_1046_),
    .B(_1057_),
    .C(_1071_),
    .D(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__nand3_2 _4383_ (.A(_1031_),
    .B(_3113_),
    .C(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__o21a_1 _4384_ (.A1(_0436_),
    .A2(_0525_),
    .B1(_2776_),
    .X(_1091_));
 sky130_fd_sc_hd__a22o_1 _4385_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(_1090_),
    .B2(_1091_),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_1 _4386_ (.A1(_2854_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .B1(_2857_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_1092_));
 sky130_fd_sc_hd__a221oi_1 _4387_ (.A1(_0589_),
    .A2(_0824_),
    .B1(_2966_),
    .B2(_0825_),
    .C1(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__nand2_1 _4388_ (.A(_2838_),
    .B(_3005_),
    .Y(_1094_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_2845_),
    .B(_0695_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _4390_ (.A(_1094_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__a221oi_2 _4391_ (.A1(_2886_),
    .A2(_2827_),
    .B1(_0537_),
    .B2(_2832_),
    .C1(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__inv_2 _4392_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1098_));
 sky130_fd_sc_hd__nand2_1 _4393_ (.A(_2879_),
    .B(_2790_),
    .Y(_1099_));
 sky130_fd_sc_hd__o221a_1 _4394_ (.A1(_2871_),
    .A2(_2870_),
    .B1(_1098_),
    .B2(_2875_),
    .C1(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__nand2_1 _4395_ (.A(_2890_),
    .B(_2777_),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2_1 _4396_ (.A(_2894_),
    .B(_2810_),
    .Y(_1102_));
 sky130_fd_sc_hd__nand2_1 _4397_ (.A(_1101_),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__a221oi_1 _4398_ (.A1(_2885_),
    .A2(_2880_),
    .B1(_2888_),
    .B2(_2802_),
    .C1(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__and4_1 _4399_ (.A(_1093_),
    .B(_1097_),
    .C(_1100_),
    .D(_1104_),
    .X(_1105_));
 sky130_fd_sc_hd__o22ai_1 _4400_ (.A1(_0796_),
    .A2(_2911_),
    .B1(_0448_),
    .B2(_2916_),
    .Y(_1106_));
 sky130_fd_sc_hd__a221oi_1 _4401_ (.A1(_3009_),
    .A2(_2903_),
    .B1(_3013_),
    .B2(_2907_),
    .C1(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__nand2_1 _4402_ (.A(_2925_),
    .B(_2806_),
    .Y(_1108_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_2928_),
    .B(_2800_),
    .Y(_1109_));
 sky130_fd_sc_hd__nand2_1 _4404_ (.A(_1108_),
    .B(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__a221oi_2 _4405_ (.A1(_2920_),
    .A2(_2891_),
    .B1(_2923_),
    .B2(_2808_),
    .C1(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_2944_),
    .B(_2798_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_1 _4407_ (.A(_2948_),
    .B(_2814_),
    .Y(_1113_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(_1112_),
    .B(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__a221oi_1 _4409_ (.A1(_0746_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2804_),
    .C1(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__nand2_1 _4410_ (.A(_2961_),
    .B(_2846_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_2965_),
    .B(_0507_),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2_1 _4412_ (.A(_1116_),
    .B(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__a221oi_1 _4413_ (.A1(_2904_),
    .A2(_2955_),
    .B1(_0334_),
    .B2(_2959_),
    .C1(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__and4_1 _4414_ (.A(_1107_),
    .B(_1111_),
    .C(_1115_),
    .D(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__nand2_1 _4415_ (.A(_2986_),
    .B(_3147_),
    .Y(_1121_));
 sky130_fd_sc_hd__o21ai_1 _4416_ (.A1(_0609_),
    .A2(_2984_),
    .B1(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__a221oi_1 _4417_ (.A1(_2908_),
    .A2(_2976_),
    .B1(_2839_),
    .B2(_2981_),
    .C1(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__or2_1 _4418_ (.A(_0564_),
    .B(_0858_),
    .X(_1124_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_2997_),
    .B(_3134_),
    .Y(_1125_));
 sky130_fd_sc_hd__nand2_1 _4420_ (.A(_3001_),
    .B(_2962_),
    .Y(_1126_));
 sky130_fd_sc_hd__o2111a_1 _4421_ (.A1(_0607_),
    .A2(_2993_),
    .B1(_1124_),
    .C1(_1125_),
    .D1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__inv_2 _4422_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .Y(_1128_));
 sky130_fd_sc_hd__o22ai_1 _4423_ (.A1(_0571_),
    .A2(_3016_),
    .B1(_1128_),
    .B2(_3022_),
    .Y(_1129_));
 sky130_fd_sc_hd__a221oi_1 _4424_ (.A1(_0326_),
    .A2(_3008_),
    .B1(_3017_),
    .B2(_3012_),
    .C1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand2_1 _4425_ (.A(_3035_),
    .B(_2817_),
    .Y(_1131_));
 sky130_fd_sc_hd__nand2_1 _4426_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_1 _4427_ (.A(_1131_),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__a221oi_1 _4428_ (.A1(_3028_),
    .A2(_0426_),
    .B1(_0550_),
    .B2(_3033_),
    .C1(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__and4_1 _4429_ (.A(_1123_),
    .B(_1127_),
    .C(_1130_),
    .D(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__nand2_1 _4430_ (.A(_3052_),
    .B(_3127_),
    .Y(_1136_));
 sky130_fd_sc_hd__nand2_1 _4431_ (.A(_3057_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1137_));
 sky130_fd_sc_hd__nand2_1 _4432_ (.A(_1136_),
    .B(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__a221oi_1 _4433_ (.A1(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0595_),
    .C1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__nand2_1 _4434_ (.A(_3069_),
    .B(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _4435_ (.A(_3072_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1141_));
 sky130_fd_sc_hd__nand2_1 _4436_ (.A(_1140_),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__a221oi_1 _4437_ (.A1(_3063_),
    .A2(_3098_),
    .B1(_3066_),
    .B2(_0352_),
    .C1(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(_3088_),
    .B(_0566_),
    .Y(_1144_));
 sky130_fd_sc_hd__o21ai_1 _4439_ (.A1(_0543_),
    .A2(_3086_),
    .B1(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__a221oi_1 _4440_ (.A1(_3077_),
    .A2(_2998_),
    .B1(_0634_),
    .B2(_3082_),
    .C1(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(_3100_),
    .B(_0707_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(_3103_),
    .B(_0649_),
    .Y(_1148_));
 sky130_fd_sc_hd__nand2_1 _4443_ (.A(_1147_),
    .B(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__a221oi_1 _4444_ (.A1(_0345_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0379_),
    .C1(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__and4_1 _4445_ (.A(_1139_),
    .B(_1143_),
    .C(_1146_),
    .D(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__and4_1 _4446_ (.A(_1105_),
    .B(_1120_),
    .C(_1135_),
    .D(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(_3126_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_1153_));
 sky130_fd_sc_hd__o21ai_1 _4448_ (.A1(_1043_),
    .A2(_3124_),
    .B1(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__a221oi_1 _4449_ (.A1(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .A2(_3117_),
    .B1(_0479_),
    .B2(_3121_),
    .C1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__or2_1 _4450_ (.A(_0880_),
    .B(_3137_),
    .X(_1156_));
 sky130_fd_sc_hd__or2_1 _4451_ (.A(_0590_),
    .B(_3141_),
    .X(_1157_));
 sky130_fd_sc_hd__nand2_1 _4452_ (.A(_3144_),
    .B(_0364_),
    .Y(_1158_));
 sky130_fd_sc_hd__o2111a_1 _4453_ (.A1(_0764_),
    .A2(_3133_),
    .B1(_1156_),
    .C1(_1157_),
    .D1(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__nand2_1 _4454_ (.A(_0325_),
    .B(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_1160_));
 sky130_fd_sc_hd__nand2_1 _4455_ (.A(_0329_),
    .B(_0459_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4456_ (.A(_1160_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__a221oi_1 _4457_ (.A1(_0384_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0422_),
    .C1(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__inv_2 _4458_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .Y(_1164_));
 sky130_fd_sc_hd__o22ai_1 _4459_ (.A1(_1164_),
    .A2(_0344_),
    .B1(_0514_),
    .B2(_0348_),
    .Y(_1165_));
 sky130_fd_sc_hd__a221oi_1 _4460_ (.A1(_0768_),
    .A2(_0337_),
    .B1(_0623_),
    .B2(_0341_),
    .C1(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__and4_1 _4461_ (.A(_1155_),
    .B(_1159_),
    .C(_1163_),
    .D(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__o22ai_1 _4462_ (.A1(_0511_),
    .A2(_0908_),
    .B1(_0815_),
    .B2(_0909_),
    .Y(_1168_));
 sky130_fd_sc_hd__a221oi_1 _4463_ (.A1(_0884_),
    .A2(_0906_),
    .B1(_0484_),
    .B2(_0907_),
    .C1(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__o22ai_1 _4464_ (.A1(_0675_),
    .A2(_0483_),
    .B1(_0921_),
    .B2(_0487_),
    .Y(_1170_));
 sky130_fd_sc_hd__a221oi_1 _4465_ (.A1(_0584_),
    .A2(_0478_),
    .B1(_3067_),
    .B2(_0480_),
    .C1(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__o22ai_1 _4466_ (.A1(_0534_),
    .A2(_0503_),
    .B1(_1060_),
    .B2(_0915_),
    .Y(_1172_));
 sky130_fd_sc_hd__a22o_1 _4467_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .B1(_0918_),
    .B2(_2792_),
    .X(_1173_));
 sky130_fd_sc_hd__nor2_1 _4468_ (.A(_1172_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__o22ai_1 _4469_ (.A1(_0676_),
    .A2(_0922_),
    .B1(_3122_),
    .B2(_0923_),
    .Y(_1175_));
 sky130_fd_sc_hd__a22o_1 _4470_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .B1(_0926_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_1176_));
 sky130_fd_sc_hd__nor2_1 _4471_ (.A(_1175_),
    .B(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__and4_1 _4472_ (.A(_1169_),
    .B(_1171_),
    .C(_1174_),
    .D(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__o22ai_1 _4473_ (.A1(_0570_),
    .A2(_0450_),
    .B1(_0655_),
    .B2(_0454_),
    .Y(_1179_));
 sky130_fd_sc_hd__a221oi_1 _4474_ (.A1(_2912_),
    .A2(_0930_),
    .B1(_0451_),
    .B2(_0931_),
    .C1(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__inv_2 _4475_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_1181_));
 sky130_fd_sc_hd__o22ai_1 _4476_ (.A1(_1181_),
    .A2(_0464_),
    .B1(_0462_),
    .B2(_0467_),
    .Y(_1182_));
 sky130_fd_sc_hd__a221oi_1 _4477_ (.A1(_3036_),
    .A2(_0936_),
    .B1(_0443_),
    .B2(_0937_),
    .C1(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _4478_ (.A(_0438_),
    .B(_0651_),
    .Y(_1184_));
 sky130_fd_sc_hd__nand2_1 _4479_ (.A(_0442_),
    .B(_2865_),
    .Y(_1185_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(_1184_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a221oi_1 _4481_ (.A1(_3083_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_0647_),
    .C1(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_0421_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1188_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(_0425_),
    .B(_0596_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _4484_ (.A(_1188_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__a221oi_1 _4485_ (.A1(_0415_),
    .A2(_0613_),
    .B1(_0418_),
    .B2(_3029_),
    .C1(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__and4_1 _4486_ (.A(_1180_),
    .B(_1183_),
    .C(_1187_),
    .D(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__nand2_1 _4487_ (.A(_0360_),
    .B(_0395_),
    .Y(_1193_));
 sky130_fd_sc_hd__nand2_1 _4488_ (.A(_0363_),
    .B(_0475_),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _4489_ (.A(_1193_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__a221oi_1 _4490_ (.A1(_0574_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0745_),
    .C1(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__nand2b_1 _4491_ (.A_N(_0369_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_1 _4492_ (.A(_0372_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1198_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(_0375_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1199_));
 sky130_fd_sc_hd__nand2_1 _4494_ (.A(_0378_),
    .B(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_1200_));
 sky130_fd_sc_hd__and4_1 _4495_ (.A(_1197_),
    .B(_1198_),
    .C(_1199_),
    .D(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__nand2_1 _4496_ (.A(_0390_),
    .B(_0385_),
    .Y(_1202_));
 sky130_fd_sc_hd__nand2_1 _4497_ (.A(_0394_),
    .B(_0416_),
    .Y(_1203_));
 sky130_fd_sc_hd__nand2_1 _4498_ (.A(_1202_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__a221oi_1 _4499_ (.A1(_0383_),
    .A2(_3092_),
    .B1(_0419_),
    .B2(_0388_),
    .C1(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__a22o_1 _4500_ (.A1(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_1206_));
 sky130_fd_sc_hd__a22o_1 _4501_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .B1(_0409_),
    .B2(_0439_),
    .X(_1207_));
 sky130_fd_sc_hd__nor2_1 _4502_ (.A(_1206_),
    .B(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__and4_1 _4503_ (.A(_1196_),
    .B(_1201_),
    .C(_1205_),
    .D(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__and4_1 _4504_ (.A(_1167_),
    .B(_1178_),
    .C(_1192_),
    .D(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__nand3_2 _4505_ (.A(_1152_),
    .B(_3113_),
    .C(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__o21a_1 _4506_ (.A1(_0648_),
    .A2(_0525_),
    .B1(_2775_),
    .X(_1212_));
 sky130_fd_sc_hd__a22o_1 _4507_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B1(_1211_),
    .B2(_1212_),
    .X(_0292_));
 sky130_fd_sc_hd__a22o_1 _4508_ (.A1(_2854_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .B1(_2857_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_1213_));
 sky130_fd_sc_hd__a221oi_1 _4509_ (.A1(_0591_),
    .A2(_0824_),
    .B1(_2891_),
    .B2(_0825_),
    .C1(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _4510_ (.A(_2838_),
    .B(_3009_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_2845_),
    .B(_2880_),
    .Y(_1216_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_1215_),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__a221oi_1 _4513_ (.A1(_2966_),
    .A2(_2827_),
    .B1(_0695_),
    .B2(_2832_),
    .C1(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__inv_2 _4514_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_1219_));
 sky130_fd_sc_hd__nand2_1 _4515_ (.A(_2879_),
    .B(_2792_),
    .Y(_1220_));
 sky130_fd_sc_hd__o221a_1 _4516_ (.A1(_0534_),
    .A2(_2870_),
    .B1(_1219_),
    .B2(_2875_),
    .C1(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_2890_),
    .B(_2786_),
    .Y(_1222_));
 sky130_fd_sc_hd__nand2_1 _4518_ (.A(_2894_),
    .B(_2812_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_1 _4519_ (.A(_1222_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__a221oi_1 _4520_ (.A1(_2885_),
    .A2(_0507_),
    .B1(_2888_),
    .B2(_2804_),
    .C1(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__and4_1 _4521_ (.A(_1214_),
    .B(_1218_),
    .C(_1221_),
    .D(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__o22ai_1 _4522_ (.A1(_0933_),
    .A2(_2911_),
    .B1(_0655_),
    .B2(_2916_),
    .Y(_1227_));
 sky130_fd_sc_hd__a221oi_1 _4523_ (.A1(_3013_),
    .A2(_2903_),
    .B1(_2956_),
    .B2(_2907_),
    .C1(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_2925_),
    .B(_2808_),
    .Y(_1229_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_2928_),
    .B(_2802_),
    .Y(_1230_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(_1229_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__a221oi_1 _4527_ (.A1(_2920_),
    .A2(_0537_),
    .B1(_2923_),
    .B2(_2810_),
    .C1(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2_1 _4528_ (.A(_2944_),
    .B(_2800_),
    .Y(_1233_));
 sky130_fd_sc_hd__nand2_1 _4529_ (.A(_2948_),
    .B(_0524_),
    .Y(_1234_));
 sky130_fd_sc_hd__nand2_1 _4530_ (.A(_1233_),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__a221oi_1 _4531_ (.A1(_0410_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2806_),
    .C1(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__nand2_1 _4532_ (.A(_2961_),
    .B(_2886_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _4533_ (.A(_2965_),
    .B(_2777_),
    .Y(_1238_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_1237_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__a221oi_1 _4535_ (.A1(_0447_),
    .A2(_2955_),
    .B1(_0384_),
    .B2(_2959_),
    .C1(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__and4_1 _4536_ (.A(_1228_),
    .B(_1232_),
    .C(_1236_),
    .D(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__nand2_1 _4537_ (.A(_2986_),
    .B(_0326_),
    .Y(_1242_));
 sky130_fd_sc_hd__o21ai_1 _4538_ (.A1(_3135_),
    .A2(_2984_),
    .B1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__a221oi_1 _4539_ (.A1(_2952_),
    .A2(_2976_),
    .B1(_2899_),
    .B2(_2981_),
    .C1(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__or2_1 _4540_ (.A(_3139_),
    .B(_0858_),
    .X(_1245_));
 sky130_fd_sc_hd__nand2_1 _4541_ (.A(_2997_),
    .B(_2971_),
    .Y(_1246_));
 sky130_fd_sc_hd__nand2_1 _4542_ (.A(_3001_),
    .B(_2817_),
    .Y(_1247_));
 sky130_fd_sc_hd__o2111a_1 _4543_ (.A1(_3084_),
    .A2(_2993_),
    .B1(_1245_),
    .C1(_1246_),
    .D1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__inv_2 _4544_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .Y(_1249_));
 sky130_fd_sc_hd__o22ai_1 _4545_ (.A1(_0725_),
    .A2(_3016_),
    .B1(_1249_),
    .B2(_3022_),
    .Y(_1250_));
 sky130_fd_sc_hd__a221oi_2 _4546_ (.A1(_3017_),
    .A2(_3008_),
    .B1(_0338_),
    .B2(_3012_),
    .C1(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__nand2_1 _4547_ (.A(_3035_),
    .B(_2865_),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_1 _4548_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1253_));
 sky130_fd_sc_hd__nand2_1 _4549_ (.A(_1252_),
    .B(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__a221oi_1 _4550_ (.A1(_3028_),
    .A2(_2932_),
    .B1(_0707_),
    .B2(_3033_),
    .C1(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__and4_1 _4551_ (.A(_1244_),
    .B(_1248_),
    .C(_1251_),
    .D(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(_3052_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1257_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_3057_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1258_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(_1257_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__a221oi_1 _4555_ (.A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0745_),
    .C1(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__nand2_1 _4556_ (.A(_3069_),
    .B(_2814_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_3072_),
    .B(_0574_),
    .Y(_1262_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_1261_),
    .B(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__a221oi_1 _4559_ (.A1(_3063_),
    .A2(_0596_),
    .B1(_3066_),
    .B2(_0622_),
    .C1(_1263_),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_3088_),
    .B(_0430_),
    .Y(_1265_));
 sky130_fd_sc_hd__o21ai_1 _4561_ (.A1(_2913_),
    .A2(_3086_),
    .B1(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__a221oi_1 _4562_ (.A1(_3077_),
    .A2(_0566_),
    .B1(_0416_),
    .B2(_3082_),
    .C1(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__nand2_1 _4563_ (.A(_3100_),
    .B(_3098_),
    .Y(_1268_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_3103_),
    .B(_3002_),
    .Y(_1269_));
 sky130_fd_sc_hd__nand2_1 _4565_ (.A(_1268_),
    .B(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__a221oi_1 _4566_ (.A1(_0510_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0631_),
    .C1(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__and4_1 _4567_ (.A(_1260_),
    .B(_1264_),
    .C(_1267_),
    .D(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__and4_1 _4568_ (.A(_1226_),
    .B(_1241_),
    .C(_1256_),
    .D(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__nand2_1 _4569_ (.A(_3126_),
    .B(_3118_),
    .Y(_1274_));
 sky130_fd_sc_hd__o21ai_1 _4570_ (.A1(_1164_),
    .A2(_3124_),
    .B1(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__a221oi_2 _4571_ (.A1(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .A2(_3117_),
    .B1(_0475_),
    .B2(_3121_),
    .C1(_1275_),
    .Y(_1276_));
 sky130_fd_sc_hd__or2_1 _4572_ (.A(_2909_),
    .B(_3137_),
    .X(_1277_));
 sky130_fd_sc_hd__or2_1 _4573_ (.A(_0741_),
    .B(_3141_),
    .X(_1278_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(_3144_),
    .B(_0391_),
    .Y(_1279_));
 sky130_fd_sc_hd__o2111a_1 _4575_ (.A1(_0902_),
    .A2(_3133_),
    .B1(_1277_),
    .C1(_1278_),
    .D1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__nand2_1 _4576_ (.A(_0325_),
    .B(_0358_),
    .Y(_1281_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_0329_),
    .B(_2977_),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2_1 _4578_ (.A(_1281_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__a221oi_1 _4579_ (.A1(_3050_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_3030_),
    .C1(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__inv_2 _4580_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_1285_));
 sky130_fd_sc_hd__o22ai_1 _4581_ (.A1(_1285_),
    .A2(_0344_),
    .B1(_0676_),
    .B2(_0348_),
    .Y(_1286_));
 sky130_fd_sc_hd__a221oi_1 _4582_ (.A1(_3092_),
    .A2(_0337_),
    .B1(_0768_),
    .B2(_0341_),
    .C1(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__and4_1 _4583_ (.A(_1276_),
    .B(_1280_),
    .C(_1284_),
    .D(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__o22ai_1 _4584_ (.A1(_0675_),
    .A2(_0908_),
    .B1(_0921_),
    .B2(_0909_),
    .Y(_1289_));
 sky130_fd_sc_hd__a221oi_1 _4585_ (.A1(_0484_),
    .A2(_0906_),
    .B1(_0345_),
    .B2(_0907_),
    .C1(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__o22ai_1 _4586_ (.A1(_0815_),
    .A2(_0483_),
    .B1(_0514_),
    .B2(_0487_),
    .Y(_1291_));
 sky130_fd_sc_hd__a221oi_1 _4587_ (.A1(_0419_),
    .A2(_0478_),
    .B1(_0584_),
    .B2(_0480_),
    .C1(_1291_),
    .Y(_1292_));
 sky130_fd_sc_hd__o22ai_1 _4588_ (.A1(_0692_),
    .A2(_0503_),
    .B1(_1181_),
    .B2(_0915_),
    .Y(_1293_));
 sky130_fd_sc_hd__a22o_1 _4589_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .B1(_0918_),
    .B2(_2794_),
    .X(_1294_));
 sky130_fd_sc_hd__nor2_1 _4590_ (.A(_1293_),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__o22ai_1 _4591_ (.A1(_0816_),
    .A2(_0922_),
    .B1(_0342_),
    .B2(_0923_),
    .Y(_1296_));
 sky130_fd_sc_hd__a22o_1 _4592_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .B1(_0926_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_1297_));
 sky130_fd_sc_hd__nor2_1 _4593_ (.A(_1296_),
    .B(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__and4_1 _4594_ (.A(_1290_),
    .B(_1292_),
    .C(_1295_),
    .D(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__o22ai_1 _4595_ (.A1(_0724_),
    .A2(_0450_),
    .B1(_0795_),
    .B2(_0454_),
    .Y(_1300_));
 sky130_fd_sc_hd__a221oi_1 _4596_ (.A1(_0451_),
    .A2(_0930_),
    .B1(_2839_),
    .B2(_0931_),
    .C1(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_2 _4597_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_1302_));
 sky130_fd_sc_hd__o22ai_1 _4598_ (.A1(_1302_),
    .A2(_0464_),
    .B1(_0660_),
    .B2(_0467_),
    .Y(_1303_));
 sky130_fd_sc_hd__a221oi_1 _4599_ (.A1(_0443_),
    .A2(_0936_),
    .B1(_0651_),
    .B2(_0937_),
    .C1(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _4600_ (.A(_0438_),
    .B(_0791_),
    .Y(_1305_));
 sky130_fd_sc_hd__nand2_1 _4601_ (.A(_0442_),
    .B(_2921_),
    .Y(_1306_));
 sky130_fd_sc_hd__nand2_1 _4602_ (.A(_1305_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__a221oi_1 _4603_ (.A1(_0457_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_0330_),
    .C1(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__nand2_1 _4604_ (.A(_0421_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1309_));
 sky130_fd_sc_hd__nand2_1 _4605_ (.A(_0425_),
    .B(_0746_),
    .Y(_1310_));
 sky130_fd_sc_hd__nand2_1 _4606_ (.A(_1309_),
    .B(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__a221oi_1 _4607_ (.A1(_0415_),
    .A2(_0352_),
    .B1(_0418_),
    .B2(_0422_),
    .C1(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__and4_1 _4608_ (.A(_1301_),
    .B(_1304_),
    .C(_1308_),
    .D(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__nand2_1 _4609_ (.A(_0360_),
    .B(_0479_),
    .Y(_1314_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(_0363_),
    .B(_0385_),
    .Y(_1315_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_1314_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__a221oi_2 _4612_ (.A1(_3064_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0884_),
    .C1(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__or2b_1 _4613_ (.A(_0368_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_1318_));
 sky130_fd_sc_hd__nand2_1 _4614_ (.A(_0371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1319_));
 sky130_fd_sc_hd__nand2_1 _4615_ (.A(_0374_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_1320_));
 sky130_fd_sc_hd__nand2_1 _4616_ (.A(_0377_),
    .B(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_1321_));
 sky130_fd_sc_hd__and4_1 _4617_ (.A(_1318_),
    .B(_1319_),
    .C(_1320_),
    .D(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__nand2_1 _4618_ (.A(_0389_),
    .B(_0634_),
    .Y(_1323_));
 sky130_fd_sc_hd__nand2_1 _4619_ (.A(_0393_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_1323_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__a221oi_1 _4621_ (.A1(_0382_),
    .A2(_0595_),
    .B1(_0323_),
    .B2(_0387_),
    .C1(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__a22o_1 _4622_ (.A1(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .A2(_0400_),
    .B1(_0403_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_1327_));
 sky130_fd_sc_hd__a22o_1 _4623_ (.A1(_0406_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .B1(_0408_),
    .B2(_0649_),
    .X(_1328_));
 sky130_fd_sc_hd__nor2_1 _4624_ (.A(_1327_),
    .B(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__and4_1 _4625_ (.A(_1317_),
    .B(_1322_),
    .C(_1326_),
    .D(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__and4_1 _4626_ (.A(_1288_),
    .B(_1299_),
    .C(_1313_),
    .D(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__nand3_2 _4627_ (.A(_1273_),
    .B(_3113_),
    .C(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__o21a_1 _4628_ (.A1(_2998_),
    .A2(_0525_),
    .B1(_2775_),
    .X(_1333_));
 sky130_fd_sc_hd__a22o_1 _4629_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B1(_1332_),
    .B2(_1333_),
    .X(_0291_));
 sky130_fd_sc_hd__a22o_1 _4630_ (.A1(_2854_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .B1(_2857_),
    .B2(_0589_),
    .X(_1334_));
 sky130_fd_sc_hd__a221oi_1 _4631_ (.A1(_0436_),
    .A2(_0824_),
    .B1(_0537_),
    .B2(_0825_),
    .C1(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_1 _4632_ (.A(_2838_),
    .B(_3013_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand2_1 _4633_ (.A(_2845_),
    .B(_0507_),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2_1 _4634_ (.A(_1336_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__a221oi_1 _4635_ (.A1(_2891_),
    .A2(_2827_),
    .B1(_2880_),
    .B2(_2832_),
    .C1(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__inv_2 _4636_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1340_));
 sky130_fd_sc_hd__nand2_1 _4637_ (.A(_2879_),
    .B(_2794_),
    .Y(_1341_));
 sky130_fd_sc_hd__o221a_1 _4638_ (.A1(_0692_),
    .A2(_2870_),
    .B1(_1340_),
    .B2(_2875_),
    .C1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__nand2_1 _4639_ (.A(_2890_),
    .B(_2788_),
    .Y(_1343_));
 sky130_fd_sc_hd__nand2_1 _4640_ (.A(_2894_),
    .B(_2814_),
    .Y(_1344_));
 sky130_fd_sc_hd__nand2_1 _4641_ (.A(_1343_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__a221oi_1 _4642_ (.A1(_2885_),
    .A2(_2777_),
    .B1(_2888_),
    .B2(_2806_),
    .C1(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__and4_1 _4643_ (.A(_1335_),
    .B(_1339_),
    .C(_1342_),
    .D(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__o22ai_1 _4644_ (.A1(_0448_),
    .A2(_2911_),
    .B1(_0795_),
    .B2(_2916_),
    .Y(_1348_));
 sky130_fd_sc_hd__a221oi_1 _4645_ (.A1(_2956_),
    .A2(_2903_),
    .B1(_3147_),
    .B2(_2907_),
    .C1(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_1 _4646_ (.A(_2925_),
    .B(_2810_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4647_ (.A(_2928_),
    .B(_2804_),
    .Y(_1351_));
 sky130_fd_sc_hd__nand2_1 _4648_ (.A(_1350_),
    .B(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__a221oi_2 _4649_ (.A1(_2920_),
    .A2(_0695_),
    .B1(_2923_),
    .B2(_2812_),
    .C1(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand2_1 _4650_ (.A(_2944_),
    .B(_2802_),
    .Y(_1354_));
 sky130_fd_sc_hd__nand2_1 _4651_ (.A(_2948_),
    .B(_3078_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_1 _4652_ (.A(_1354_),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__a221oi_1 _4653_ (.A1(_3104_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2808_),
    .C1(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__nand2_1 _4654_ (.A(_2961_),
    .B(_2966_),
    .Y(_1358_));
 sky130_fd_sc_hd__nand2_1 _4655_ (.A(_2965_),
    .B(_2786_),
    .Y(_1359_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_1358_),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__a221oi_1 _4657_ (.A1(_2987_),
    .A2(_2955_),
    .B1(_3050_),
    .B2(_2959_),
    .C1(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__and4_1 _4658_ (.A(_1349_),
    .B(_1353_),
    .C(_1357_),
    .D(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__nand2_1 _4659_ (.A(_2986_),
    .B(_3017_),
    .Y(_1363_));
 sky130_fd_sc_hd__o21ai_1 _4660_ (.A1(_0607_),
    .A2(_2984_),
    .B1(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__a221oi_1 _4661_ (.A1(_2912_),
    .A2(_2976_),
    .B1(_2904_),
    .B2(_2981_),
    .C1(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__or2_1 _4662_ (.A(_0609_),
    .B(_0858_),
    .X(_1366_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_2997_),
    .B(_3083_),
    .Y(_1367_));
 sky130_fd_sc_hd__nand2_1 _4664_ (.A(_3001_),
    .B(_2865_),
    .Y(_1368_));
 sky130_fd_sc_hd__o2111a_1 _4665_ (.A1(_0590_),
    .A2(_2993_),
    .B1(_1366_),
    .C1(_1367_),
    .D1(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__inv_2 _4666_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_1370_));
 sky130_fd_sc_hd__o22ai_1 _4667_ (.A1(_0864_),
    .A2(_3016_),
    .B1(_1370_),
    .B2(_3022_),
    .Y(_1371_));
 sky130_fd_sc_hd__a221oi_1 _4668_ (.A1(_0338_),
    .A2(_3008_),
    .B1(_0334_),
    .B2(_3012_),
    .C1(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_1 _4669_ (.A(_3035_),
    .B(_2921_),
    .Y(_1373_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1374_));
 sky130_fd_sc_hd__nand2_1 _4671_ (.A(_1373_),
    .B(_1374_),
    .Y(_1375_));
 sky130_fd_sc_hd__a221oi_1 _4672_ (.A1(_3028_),
    .A2(_0550_),
    .B1(_3098_),
    .B2(_3033_),
    .C1(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__and4_1 _4673_ (.A(_1365_),
    .B(_1369_),
    .C(_1372_),
    .D(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_3052_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _4675_ (.A(_3057_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_1 _4676_ (.A(_1378_),
    .B(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__a221oi_2 _4677_ (.A1(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0884_),
    .C1(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _4678_ (.A(_3069_),
    .B(_0524_),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _4679_ (.A(_3072_),
    .B(_3064_),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_1 _4680_ (.A(_1382_),
    .B(_1383_),
    .Y(_1384_));
 sky130_fd_sc_hd__a221oi_1 _4681_ (.A1(_3063_),
    .A2(_0746_),
    .B1(_3066_),
    .B2(_3029_),
    .C1(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _4682_ (.A(_3088_),
    .B(_0647_),
    .Y(_1386_));
 sky130_fd_sc_hd__o21ai_1 _4683_ (.A1(_0452_),
    .A2(_3086_),
    .B1(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__a221oi_1 _4684_ (.A1(_3077_),
    .A2(_0430_),
    .B1(_3067_),
    .B2(_3082_),
    .C1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__nand2_1 _4685_ (.A(_3100_),
    .B(_0596_),
    .Y(_1389_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(_3103_),
    .B(_3036_),
    .Y(_1390_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_1389_),
    .B(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a221oi_1 _4688_ (.A1(_3053_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0471_),
    .C1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__and4_2 _4689_ (.A(_1381_),
    .B(_1385_),
    .C(_1388_),
    .D(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__and4_1 _4690_ (.A(_1347_),
    .B(_1362_),
    .C(_1377_),
    .D(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__nand2_1 _4691_ (.A(_3126_),
    .B(_0364_),
    .Y(_1395_));
 sky130_fd_sc_hd__o21ai_1 _4692_ (.A1(_1285_),
    .A2(_3124_),
    .B1(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__a221oi_1 _4693_ (.A1(_3118_),
    .A2(_3117_),
    .B1(_0385_),
    .B2(_3121_),
    .C1(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__or2_1 _4694_ (.A(_0543_),
    .B(_3137_),
    .X(_1398_));
 sky130_fd_sc_hd__or2_1 _4695_ (.A(_0880_),
    .B(_3141_),
    .X(_1399_));
 sky130_fd_sc_hd__nand2_1 _4696_ (.A(_3144_),
    .B(_3079_),
    .Y(_1400_));
 sky130_fd_sc_hd__o2111a_1 _4697_ (.A1(_1043_),
    .A2(_3133_),
    .B1(_1398_),
    .C1(_1399_),
    .D1(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__nand2_1 _4698_ (.A(_0325_),
    .B(_0623_),
    .Y(_1402_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(_0329_),
    .B(_2908_),
    .Y(_1403_));
 sky130_fd_sc_hd__nand2_1 _4700_ (.A(_1402_),
    .B(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__a221oi_1 _4701_ (.A1(_0358_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0574_),
    .C1(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__inv_2 _4702_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_1406_));
 sky130_fd_sc_hd__o22ai_1 _4703_ (.A1(_1406_),
    .A2(_0344_),
    .B1(_0816_),
    .B2(_0348_),
    .Y(_1407_));
 sky130_fd_sc_hd__a221oi_1 _4704_ (.A1(_0595_),
    .A2(_0337_),
    .B1(_3092_),
    .B2(_0341_),
    .C1(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__and4_1 _4705_ (.A(_1397_),
    .B(_1401_),
    .C(_1405_),
    .D(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__o22ai_1 _4706_ (.A1(_0815_),
    .A2(_0908_),
    .B1(_0514_),
    .B2(_0909_),
    .Y(_1410_));
 sky130_fd_sc_hd__a221oi_1 _4707_ (.A1(_0345_),
    .A2(_0906_),
    .B1(_0510_),
    .B2(_0907_),
    .C1(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__o22ai_1 _4708_ (.A1(_0921_),
    .A2(_0483_),
    .B1(_0676_),
    .B2(_0487_),
    .Y(_1412_));
 sky130_fd_sc_hd__a221oi_1 _4709_ (.A1(_0323_),
    .A2(_0478_),
    .B1(_0419_),
    .B2(_0480_),
    .C1(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__o22ai_1 _4710_ (.A1(_0832_),
    .A2(_0503_),
    .B1(_1302_),
    .B2(_0915_),
    .Y(_1414_));
 sky130_fd_sc_hd__a22o_1 _4711_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .B1(_0918_),
    .B2(_2796_),
    .X(_1415_));
 sky130_fd_sc_hd__nor2_1 _4712_ (.A(_1414_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__o22ai_1 _4713_ (.A1(_3131_),
    .A2(_0922_),
    .B1(_0618_),
    .B2(_0923_),
    .Y(_1417_));
 sky130_fd_sc_hd__a22o_1 _4714_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .B1(_0926_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_1418_));
 sky130_fd_sc_hd__nor2_1 _4715_ (.A(_1417_),
    .B(_1418_),
    .Y(_1419_));
 sky130_fd_sc_hd__and4_1 _4716_ (.A(_1411_),
    .B(_1413_),
    .C(_1416_),
    .D(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__o22ai_1 _4717_ (.A1(_0863_),
    .A2(_0450_),
    .B1(_0932_),
    .B2(_0454_),
    .Y(_1421_));
 sky130_fd_sc_hd__a221oi_1 _4718_ (.A1(_2839_),
    .A2(_0930_),
    .B1(_2899_),
    .B2(_0931_),
    .C1(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_1423_));
 sky130_fd_sc_hd__o22ai_1 _4720_ (.A1(_1423_),
    .A2(_0464_),
    .B1(_0800_),
    .B2(_0467_),
    .Y(_1424_));
 sky130_fd_sc_hd__a221oi_1 _4721_ (.A1(_0651_),
    .A2(_0936_),
    .B1(_0791_),
    .B2(_0937_),
    .C1(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__nand2_1 _4722_ (.A(_0438_),
    .B(_2962_),
    .Y(_1426_));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(_0442_),
    .B(_2828_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_1 _4724_ (.A(_1426_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__a221oi_1 _4725_ (.A1(_0459_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_3134_),
    .C1(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__nand2_1 _4726_ (.A(_0421_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_1 _4727_ (.A(_0425_),
    .B(_0410_),
    .Y(_1431_));
 sky130_fd_sc_hd__nand2_1 _4728_ (.A(_1430_),
    .B(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__a221oi_1 _4729_ (.A1(_0415_),
    .A2(_0622_),
    .B1(_0418_),
    .B2(_3030_),
    .C1(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__and4_1 _4730_ (.A(_1422_),
    .B(_1425_),
    .C(_1429_),
    .D(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(_0360_),
    .B(_0475_),
    .Y(_1435_));
 sky130_fd_sc_hd__nand2_1 _4732_ (.A(_0363_),
    .B(_0634_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_1435_),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__a221oi_1 _4734_ (.A1(_0426_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0484_),
    .C1(_1437_),
    .Y(_1438_));
 sky130_fd_sc_hd__or2b_1 _4735_ (.A(_0368_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_1439_));
 sky130_fd_sc_hd__nand2_1 _4736_ (.A(_0371_),
    .B(_0379_),
    .Y(_1440_));
 sky130_fd_sc_hd__nand2_1 _4737_ (.A(_0374_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_1441_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0377_),
    .B(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_1442_));
 sky130_fd_sc_hd__and4_1 _4739_ (.A(_1439_),
    .B(_1440_),
    .C(_1441_),
    .D(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__nand2_1 _4740_ (.A(_0389_),
    .B(_0416_),
    .Y(_1444_));
 sky130_fd_sc_hd__nand2_1 _4741_ (.A(_0393_),
    .B(_0584_),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _4742_ (.A(_1444_),
    .B(_1445_),
    .Y(_1446_));
 sky130_fd_sc_hd__a221oi_1 _4743_ (.A1(_0382_),
    .A2(_0745_),
    .B1(_0613_),
    .B2(_0387_),
    .C1(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__a22o_1 _4744_ (.A1(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .A2(_0400_),
    .B1(_0403_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_1448_));
 sky130_fd_sc_hd__a22o_1 _4745_ (.A1(_0406_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .B1(_0408_),
    .B2(_3002_),
    .X(_1449_));
 sky130_fd_sc_hd__nor2_1 _4746_ (.A(_1448_),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__and4_1 _4747_ (.A(_1438_),
    .B(_1443_),
    .C(_1447_),
    .D(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__and4_1 _4748_ (.A(_1409_),
    .B(_1420_),
    .C(_1434_),
    .D(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__nand3_2 _4749_ (.A(_1394_),
    .B(_3113_),
    .C(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__o21a_1 _4750_ (.A1(_0566_),
    .A2(_3112_),
    .B1(_2775_),
    .X(_1454_));
 sky130_fd_sc_hd__a22o_1 _4751_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B1(_1453_),
    .B2(_1454_),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_1 _4752_ (.A1(_2854_),
    .A2(_0436_),
    .B1(_2857_),
    .B2(_0591_),
    .X(_1455_));
 sky130_fd_sc_hd__a221oi_1 _4753_ (.A1(_0648_),
    .A2(_0824_),
    .B1(_0695_),
    .B2(_0825_),
    .C1(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__nand2_1 _4754_ (.A(_2838_),
    .B(_2956_),
    .Y(_1457_));
 sky130_fd_sc_hd__nand2_1 _4755_ (.A(_2845_),
    .B(_2777_),
    .Y(_1458_));
 sky130_fd_sc_hd__nand2_1 _4756_ (.A(_1457_),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__a221oi_1 _4757_ (.A1(_0537_),
    .A2(_2827_),
    .B1(_0507_),
    .B2(_2832_),
    .C1(_1459_),
    .Y(_1460_));
 sky130_fd_sc_hd__inv_2 _4758_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1461_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(_2879_),
    .B(_2796_),
    .Y(_1462_));
 sky130_fd_sc_hd__o221a_1 _4760_ (.A1(_0832_),
    .A2(_2870_),
    .B1(_1461_),
    .B2(_2875_),
    .C1(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__nand2_1 _4761_ (.A(_2890_),
    .B(_2790_),
    .Y(_1464_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(_2894_),
    .B(_0524_),
    .Y(_1465_));
 sky130_fd_sc_hd__nand2_1 _4763_ (.A(_1464_),
    .B(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__a221oi_1 _4764_ (.A1(_2885_),
    .A2(_2786_),
    .B1(_2888_),
    .B2(_2808_),
    .C1(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__and4_1 _4765_ (.A(_1456_),
    .B(_1460_),
    .C(_1463_),
    .D(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__o22ai_1 _4766_ (.A1(_0655_),
    .A2(_2911_),
    .B1(_0932_),
    .B2(_2916_),
    .Y(_1469_));
 sky130_fd_sc_hd__a221oi_1 _4767_ (.A1(_3147_),
    .A2(_2903_),
    .B1(_0326_),
    .B2(_2907_),
    .C1(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_2925_),
    .B(_2812_),
    .Y(_1471_));
 sky130_fd_sc_hd__nand2_1 _4769_ (.A(_2928_),
    .B(_2806_),
    .Y(_1472_));
 sky130_fd_sc_hd__nand2_1 _4770_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__a221oi_1 _4771_ (.A1(_2920_),
    .A2(_2880_),
    .B1(_2923_),
    .B2(_2814_),
    .C1(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _4772_ (.A(_2944_),
    .B(_2804_),
    .Y(_1475_));
 sky130_fd_sc_hd__nand2_1 _4773_ (.A(_2948_),
    .B(_0589_),
    .Y(_1476_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_1475_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__a221oi_1 _4775_ (.A1(_0379_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2810_),
    .C1(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__nand2_1 _4776_ (.A(_2961_),
    .B(_2891_),
    .Y(_1479_));
 sky130_fd_sc_hd__nand2_1 _4777_ (.A(_2965_),
    .B(_2788_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2_1 _4778_ (.A(_1479_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__a221oi_1 _4779_ (.A1(_3005_),
    .A2(_2955_),
    .B1(_0358_),
    .B2(_2959_),
    .C1(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__and4_1 _4780_ (.A(_1470_),
    .B(_1474_),
    .C(_1478_),
    .D(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_2986_),
    .B(_0338_),
    .Y(_1484_));
 sky130_fd_sc_hd__o21ai_1 _4782_ (.A1(_3084_),
    .A2(_2984_),
    .B1(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__a221oi_1 _4783_ (.A1(_0451_),
    .A2(_2976_),
    .B1(_0447_),
    .B2(_2981_),
    .C1(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__or2_1 _4784_ (.A(_3135_),
    .B(_0858_),
    .X(_1487_));
 sky130_fd_sc_hd__nand2_1 _4785_ (.A(_2997_),
    .B(_0457_),
    .Y(_1488_));
 sky130_fd_sc_hd__nand2_1 _4786_ (.A(_3001_),
    .B(_2921_),
    .Y(_1489_));
 sky130_fd_sc_hd__o2111a_1 _4787_ (.A1(_0741_),
    .A2(_2993_),
    .B1(_1487_),
    .C1(_1488_),
    .D1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__inv_2 _4788_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_1491_));
 sky130_fd_sc_hd__o22ai_1 _4789_ (.A1(_1007_),
    .A2(_3016_),
    .B1(_1491_),
    .B2(_3022_),
    .Y(_1492_));
 sky130_fd_sc_hd__a221oi_1 _4790_ (.A1(_0334_),
    .A2(_3008_),
    .B1(_0384_),
    .B2(_3012_),
    .C1(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__nand2_1 _4791_ (.A(_3035_),
    .B(_2828_),
    .Y(_1494_));
 sky130_fd_sc_hd__nand2_1 _4792_ (.A(_3039_),
    .B(_0550_),
    .Y(_1495_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_1494_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__a221oi_1 _4794_ (.A1(_3028_),
    .A2(_0707_),
    .B1(_0596_),
    .B2(_3033_),
    .C1(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__and4_1 _4795_ (.A(_1486_),
    .B(_1490_),
    .C(_1493_),
    .D(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__nand2_1 _4796_ (.A(_3052_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1499_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(_3057_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_1500_));
 sky130_fd_sc_hd__nand2_1 _4798_ (.A(_1499_),
    .B(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__a221oi_2 _4799_ (.A1(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0484_),
    .C1(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__nand2_1 _4800_ (.A(_3069_),
    .B(_3078_),
    .Y(_1503_));
 sky130_fd_sc_hd__nand2_1 _4801_ (.A(_3072_),
    .B(_0426_),
    .Y(_1504_));
 sky130_fd_sc_hd__nand2_1 _4802_ (.A(_1503_),
    .B(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__a221oi_1 _4803_ (.A1(_3063_),
    .A2(_0410_),
    .B1(_3066_),
    .B2(_0422_),
    .C1(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__nand2_1 _4804_ (.A(_3088_),
    .B(_0330_),
    .Y(_1507_));
 sky130_fd_sc_hd__o21ai_1 _4805_ (.A1(_0656_),
    .A2(_3086_),
    .B1(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__a221oi_1 _4806_ (.A1(_3077_),
    .A2(_0647_),
    .B1(_0584_),
    .B2(_3082_),
    .C1(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(_3100_),
    .B(_0746_),
    .Y(_1510_));
 sky130_fd_sc_hd__nand2_1 _4808_ (.A(_3103_),
    .B(_0443_),
    .Y(_1511_));
 sky130_fd_sc_hd__nand2_1 _4809_ (.A(_1510_),
    .B(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__a221oi_1 _4810_ (.A1(_3044_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0439_),
    .C1(_1512_),
    .Y(_1513_));
 sky130_fd_sc_hd__and4_1 _4811_ (.A(_1502_),
    .B(_1506_),
    .C(_1509_),
    .D(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__and4_2 _4812_ (.A(_1468_),
    .B(_1483_),
    .C(_1498_),
    .D(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__nand2_1 _4813_ (.A(_3126_),
    .B(_0391_),
    .Y(_1516_));
 sky130_fd_sc_hd__o21ai_1 _4814_ (.A1(_1406_),
    .A2(_3124_),
    .B1(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__a221oi_2 _4815_ (.A1(_0364_),
    .A2(_3117_),
    .B1(_0634_),
    .B2(_3121_),
    .C1(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__or2_1 _4816_ (.A(_2913_),
    .B(_3137_),
    .X(_1519_));
 sky130_fd_sc_hd__or2_1 _4817_ (.A(_2909_),
    .B(_3141_),
    .X(_1520_));
 sky130_fd_sc_hd__nand2_1 _4818_ (.A(_3144_),
    .B(_0395_),
    .Y(_1521_));
 sky130_fd_sc_hd__o2111a_1 _4819_ (.A1(_1164_),
    .A2(_3133_),
    .B1(_1519_),
    .C1(_1520_),
    .D1(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__nand2_1 _4820_ (.A(_0325_),
    .B(_0768_),
    .Y(_1523_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(_0329_),
    .B(_2952_),
    .Y(_1524_));
 sky130_fd_sc_hd__nand2_1 _4822_ (.A(_1523_),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__a221oi_1 _4823_ (.A1(_0623_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_3064_),
    .C1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__inv_2 _4824_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_1527_));
 sky130_fd_sc_hd__o22ai_1 _4825_ (.A1(_1527_),
    .A2(_0344_),
    .B1(_3131_),
    .B2(_0348_),
    .Y(_1528_));
 sky130_fd_sc_hd__a221oi_1 _4826_ (.A1(_0745_),
    .A2(_0337_),
    .B1(_0595_),
    .B2(_0341_),
    .C1(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__and4_1 _4827_ (.A(_1518_),
    .B(_1522_),
    .C(_1526_),
    .D(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__o22ai_1 _4828_ (.A1(_0921_),
    .A2(_0908_),
    .B1(_0676_),
    .B2(_0909_),
    .Y(_1531_));
 sky130_fd_sc_hd__a221oi_1 _4829_ (.A1(_0510_),
    .A2(_0906_),
    .B1(_3053_),
    .B2(_0907_),
    .C1(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__o22ai_1 _4830_ (.A1(_0514_),
    .A2(_0483_),
    .B1(_0816_),
    .B2(_0487_),
    .Y(_1533_));
 sky130_fd_sc_hd__a221oi_1 _4831_ (.A1(_0613_),
    .A2(_0478_),
    .B1(_0323_),
    .B2(_0480_),
    .C1(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__o22ai_1 _4832_ (.A1(_0977_),
    .A2(_0503_),
    .B1(_1423_),
    .B2(_0915_),
    .Y(_1535_));
 sky130_fd_sc_hd__a22o_1 _4833_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .B1(_0918_),
    .B2(_2798_),
    .X(_1536_));
 sky130_fd_sc_hd__nor2_1 _4834_ (.A(_1535_),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__o22ai_1 _4835_ (.A1(_0606_),
    .A2(_0922_),
    .B1(_0764_),
    .B2(_0923_),
    .Y(_1538_));
 sky130_fd_sc_hd__a22o_1 _4836_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .B1(_0926_),
    .B2(_0566_),
    .X(_1539_));
 sky130_fd_sc_hd__nor2_1 _4837_ (.A(_1538_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__and4_1 _4838_ (.A(_1532_),
    .B(_1534_),
    .C(_1537_),
    .D(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_0372_),
    .B(_0631_),
    .Y(_1542_));
 sky130_fd_sc_hd__o21ai_1 _4840_ (.A1(_0465_),
    .A2(_0369_),
    .B1(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__a221oi_2 _4841_ (.A1(_0651_),
    .A2(_0378_),
    .B1(_0471_),
    .B2(_0375_),
    .C1(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__nand2_1 _4842_ (.A(_0360_),
    .B(_0385_),
    .Y(_1545_));
 sky130_fd_sc_hd__nand2_1 _4843_ (.A(_0363_),
    .B(_0416_),
    .Y(_1546_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(_1545_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__a221oi_2 _4845_ (.A1(_2932_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0345_),
    .C1(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__a22o_1 _4846_ (.A1(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_1549_));
 sky130_fd_sc_hd__a22o_1 _4847_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .B1(_0409_),
    .B2(_3036_),
    .X(_1550_));
 sky130_fd_sc_hd__nor2_1 _4848_ (.A(_1549_),
    .B(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(_0390_),
    .B(_3067_),
    .Y(_1552_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1553_));
 sky130_fd_sc_hd__nand2_1 _4851_ (.A(_1552_),
    .B(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__a221oi_1 _4852_ (.A1(_0383_),
    .A2(_0884_),
    .B1(_0352_),
    .B2(_0388_),
    .C1(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__and4_1 _4853_ (.A(_1544_),
    .B(_1548_),
    .C(_1551_),
    .D(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__o22ai_1 _4854_ (.A1(_3018_),
    .A2(_0450_),
    .B1(_3014_),
    .B2(_0454_),
    .Y(_1557_));
 sky130_fd_sc_hd__a221oi_1 _4855_ (.A1(_2899_),
    .A2(_0930_),
    .B1(_2904_),
    .B2(_0931_),
    .C1(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__inv_2 _4856_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1559_));
 sky130_fd_sc_hd__o22ai_1 _4857_ (.A1(_1559_),
    .A2(_0464_),
    .B1(_0938_),
    .B2(_0467_),
    .Y(_1560_));
 sky130_fd_sc_hd__a221oi_1 _4858_ (.A1(_0791_),
    .A2(_0936_),
    .B1(_2962_),
    .B2(_0937_),
    .C1(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__nand2_1 _4859_ (.A(_0438_),
    .B(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_1562_));
 sky130_fd_sc_hd__nand2_1 _4860_ (.A(_0442_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_1563_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(_1562_),
    .B(_1563_),
    .Y(_1564_));
 sky130_fd_sc_hd__a221oi_1 _4862_ (.A1(_2977_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_2971_),
    .C1(_1564_),
    .Y(_1565_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_0421_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_1566_));
 sky130_fd_sc_hd__nand2_1 _4864_ (.A(_0425_),
    .B(_3104_),
    .Y(_1567_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(_1566_),
    .B(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__a221oi_1 _4866_ (.A1(_0415_),
    .A2(_3029_),
    .B1(_0418_),
    .B2(_0574_),
    .C1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__and4_1 _4867_ (.A(_1558_),
    .B(_1561_),
    .C(_1565_),
    .D(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__and4_1 _4868_ (.A(_1530_),
    .B(_1541_),
    .C(_1556_),
    .D(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__nand3_2 _4869_ (.A(_1515_),
    .B(_3113_),
    .C(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__o21a_1 _4870_ (.A1(_0430_),
    .A2(_3112_),
    .B1(_2775_),
    .X(_1573_));
 sky130_fd_sc_hd__a22o_1 _4871_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B1(_1572_),
    .B2(_1573_),
    .X(_0289_));
 sky130_fd_sc_hd__a22o_1 _4872_ (.A1(_2854_),
    .A2(_0648_),
    .B1(_2857_),
    .B2(_0436_),
    .X(_1574_));
 sky130_fd_sc_hd__a221oi_1 _4873_ (.A1(_2998_),
    .A2(_0824_),
    .B1(_2880_),
    .B2(_0825_),
    .C1(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__nand2_1 _4874_ (.A(_2838_),
    .B(_3147_),
    .Y(_1576_));
 sky130_fd_sc_hd__nand2_1 _4875_ (.A(_2845_),
    .B(_2786_),
    .Y(_1577_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(_1576_),
    .B(_1577_),
    .Y(_1578_));
 sky130_fd_sc_hd__a221oi_1 _4877_ (.A1(_0695_),
    .A2(_2827_),
    .B1(_2777_),
    .B2(_2832_),
    .C1(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__inv_2 _4878_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1580_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(_2879_),
    .B(_2798_),
    .Y(_1581_));
 sky130_fd_sc_hd__o221a_1 _4880_ (.A1(_0977_),
    .A2(_2869_),
    .B1(_1580_),
    .B2(_2875_),
    .C1(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__nand2_1 _4881_ (.A(_2890_),
    .B(_2792_),
    .Y(_1583_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(_2894_),
    .B(_3078_),
    .Y(_1584_));
 sky130_fd_sc_hd__nand2_1 _4883_ (.A(_1583_),
    .B(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__a221oi_1 _4884_ (.A1(_2885_),
    .A2(_2788_),
    .B1(_2888_),
    .B2(_2810_),
    .C1(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__and4_1 _4885_ (.A(_1575_),
    .B(_1579_),
    .C(_1582_),
    .D(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__o22ai_1 _4886_ (.A1(_0795_),
    .A2(_2911_),
    .B1(_3014_),
    .B2(_2916_),
    .Y(_1588_));
 sky130_fd_sc_hd__a221oi_1 _4887_ (.A1(_0326_),
    .A2(_2903_),
    .B1(_3017_),
    .B2(_2907_),
    .C1(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__nand2_1 _4888_ (.A(_2925_),
    .B(_2814_),
    .Y(_1590_));
 sky130_fd_sc_hd__nand2_1 _4889_ (.A(_2928_),
    .B(_2808_),
    .Y(_1591_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(_1590_),
    .B(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__a221oi_1 _4891_ (.A1(_2920_),
    .A2(_0507_),
    .B1(_2923_),
    .B2(_0524_),
    .C1(_1592_),
    .Y(_1593_));
 sky130_fd_sc_hd__nand2_1 _4892_ (.A(_2944_),
    .B(_2806_),
    .Y(_1594_));
 sky130_fd_sc_hd__nand2_1 _4893_ (.A(_2948_),
    .B(_0591_),
    .Y(_1595_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(_1594_),
    .B(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__a221oi_1 _4895_ (.A1(_0631_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_2812_),
    .C1(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _4896_ (.A(_2961_),
    .B(_0537_),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_1 _4897_ (.A(_2965_),
    .B(_2790_),
    .Y(_1599_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_1598_),
    .B(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__a221oi_1 _4899_ (.A1(_3009_),
    .A2(_2955_),
    .B1(_0623_),
    .B2(_2959_),
    .C1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__and4_1 _4900_ (.A(_1589_),
    .B(_1593_),
    .C(_1597_),
    .D(_1601_),
    .X(_1602_));
 sky130_fd_sc_hd__nand2_1 _4901_ (.A(_2986_),
    .B(_0334_),
    .Y(_1603_));
 sky130_fd_sc_hd__o21ai_1 _4902_ (.A1(_0590_),
    .A2(_2984_),
    .B1(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__a221oi_1 _4903_ (.A1(_2839_),
    .A2(_2976_),
    .B1(_2987_),
    .B2(_2981_),
    .C1(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__or2_1 _4904_ (.A(_0607_),
    .B(_0858_),
    .X(_1606_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_2997_),
    .B(_0459_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(_3001_),
    .B(_2828_),
    .Y(_1608_));
 sky130_fd_sc_hd__o2111a_1 _4907_ (.A1(_0880_),
    .A2(_2993_),
    .B1(_1606_),
    .C1(_1607_),
    .D1(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__o22ai_1 _4908_ (.A1(_1128_),
    .A2(_3016_),
    .B1(_0490_),
    .B2(_3022_),
    .Y(_1610_));
 sky130_fd_sc_hd__a221oi_1 _4909_ (.A1(_0384_),
    .A2(_3008_),
    .B1(_3050_),
    .B2(_3012_),
    .C1(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(_3035_),
    .B(_2846_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _4911_ (.A(_3039_),
    .B(_0707_),
    .Y(_1613_));
 sky130_fd_sc_hd__nand2_1 _4912_ (.A(_1612_),
    .B(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__a221oi_1 _4913_ (.A1(_3028_),
    .A2(_3098_),
    .B1(_0746_),
    .B2(_3033_),
    .C1(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__and4_1 _4914_ (.A(_1605_),
    .B(_1609_),
    .C(_1611_),
    .D(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__nand2_1 _4915_ (.A(_3052_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1617_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(_3057_),
    .B(_3118_),
    .Y(_1618_));
 sky130_fd_sc_hd__nand2_1 _4917_ (.A(_1617_),
    .B(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__a221oi_2 _4918_ (.A1(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0345_),
    .C1(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__nand2_1 _4919_ (.A(_3069_),
    .B(_0589_),
    .Y(_1621_));
 sky130_fd_sc_hd__nand2_1 _4920_ (.A(_3072_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1622_));
 sky130_fd_sc_hd__nand2_1 _4921_ (.A(_1621_),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__a221oi_1 _4922_ (.A1(_3063_),
    .A2(_3104_),
    .B1(_3066_),
    .B2(_3030_),
    .C1(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__nand2_1 _4923_ (.A(_3088_),
    .B(_3134_),
    .Y(_1625_));
 sky130_fd_sc_hd__o21ai_1 _4924_ (.A1(_0796_),
    .A2(_3086_),
    .B1(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__a221oi_1 _4925_ (.A1(_3077_),
    .A2(_0330_),
    .B1(_0419_),
    .B2(_3082_),
    .C1(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__nand2_1 _4926_ (.A(_3100_),
    .B(_0410_),
    .Y(_1628_));
 sky130_fd_sc_hd__nand2_1 _4927_ (.A(_3103_),
    .B(_0651_),
    .Y(_1629_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_1628_),
    .B(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__a221oi_1 _4929_ (.A1(_3058_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0649_),
    .C1(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__and4_1 _4930_ (.A(_1620_),
    .B(_1624_),
    .C(_1627_),
    .D(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__and4_1 _4931_ (.A(_1587_),
    .B(_1602_),
    .C(_1616_),
    .D(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_3126_),
    .B(_3079_),
    .Y(_1634_));
 sky130_fd_sc_hd__o21ai_1 _4933_ (.A1(_1527_),
    .A2(_3124_),
    .B1(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__a221oi_1 _4934_ (.A1(_0391_),
    .A2(_3117_),
    .B1(_0416_),
    .B2(_3121_),
    .C1(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__or2_1 _4935_ (.A(_0452_),
    .B(_3137_),
    .X(_1637_));
 sky130_fd_sc_hd__or2_1 _4936_ (.A(_0543_),
    .B(_3141_),
    .X(_1638_));
 sky130_fd_sc_hd__nand2_1 _4937_ (.A(_3144_),
    .B(_0479_),
    .Y(_1639_));
 sky130_fd_sc_hd__o2111a_1 _4938_ (.A1(_1285_),
    .A2(_3133_),
    .B1(_1637_),
    .C1(_1638_),
    .D1(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__nand2_1 _4939_ (.A(_0325_),
    .B(_3092_),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_0329_),
    .B(_2912_),
    .Y(_1642_));
 sky130_fd_sc_hd__nand2_1 _4941_ (.A(_1641_),
    .B(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__a221oi_2 _4942_ (.A1(_0768_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0426_),
    .C1(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__inv_2 _4943_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_1645_));
 sky130_fd_sc_hd__o22ai_1 _4944_ (.A1(_1645_),
    .A2(_0344_),
    .B1(_0606_),
    .B2(_0348_),
    .Y(_1646_));
 sky130_fd_sc_hd__a221oi_1 _4945_ (.A1(_0884_),
    .A2(_0337_),
    .B1(_0745_),
    .B2(_0341_),
    .C1(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__and4_1 _4946_ (.A(_1636_),
    .B(_1640_),
    .C(_1644_),
    .D(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__o22ai_1 _4947_ (.A1(_0514_),
    .A2(_0908_),
    .B1(_0816_),
    .B2(_0909_),
    .Y(_1649_));
 sky130_fd_sc_hd__a221oi_1 _4948_ (.A1(_3053_),
    .A2(_0906_),
    .B1(_3044_),
    .B2(_0907_),
    .C1(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__o22ai_1 _4949_ (.A1(_0676_),
    .A2(_0483_),
    .B1(_3131_),
    .B2(_0487_),
    .Y(_1651_));
 sky130_fd_sc_hd__a221oi_1 _4950_ (.A1(_0352_),
    .A2(_0478_),
    .B1(_0613_),
    .B2(_0480_),
    .C1(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__o22ai_1 _4951_ (.A1(_1098_),
    .A2(_0503_),
    .B1(_1559_),
    .B2(_0915_),
    .Y(_1653_));
 sky130_fd_sc_hd__a22o_1 _4952_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .B1(_0918_),
    .B2(_2800_),
    .X(_1654_));
 sky130_fd_sc_hd__nor2_1 _4953_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__o22ai_1 _4954_ (.A1(_3122_),
    .A2(_0922_),
    .B1(_0902_),
    .B2(_0923_),
    .Y(_1656_));
 sky130_fd_sc_hd__a22o_1 _4955_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .B1(_0926_),
    .B2(_0430_),
    .X(_1657_));
 sky130_fd_sc_hd__nor2_1 _4956_ (.A(_1656_),
    .B(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__and4_1 _4957_ (.A(_1650_),
    .B(_1652_),
    .C(_1655_),
    .D(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__nand2_1 _4958_ (.A(_0372_),
    .B(_0471_),
    .Y(_1660_));
 sky130_fd_sc_hd__o21ai_1 _4959_ (.A1(_0661_),
    .A2(_0369_),
    .B1(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__a221oi_1 _4960_ (.A1(_0791_),
    .A2(_0378_),
    .B1(_0439_),
    .B2(_0375_),
    .C1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__nand2_1 _4961_ (.A(_0360_),
    .B(_0634_),
    .Y(_1663_));
 sky130_fd_sc_hd__nand2_1 _4962_ (.A(_0363_),
    .B(_3067_),
    .Y(_1664_));
 sky130_fd_sc_hd__nand2_1 _4963_ (.A(_1663_),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__a221oi_1 _4964_ (.A1(_0550_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0510_),
    .C1(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__a22o_1 _4965_ (.A1(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_1667_));
 sky130_fd_sc_hd__a22o_1 _4966_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .B1(_0409_),
    .B2(_0443_),
    .X(_1668_));
 sky130_fd_sc_hd__nor2_1 _4967_ (.A(_1667_),
    .B(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(_0390_),
    .B(_0584_),
    .Y(_1670_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_1671_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_1670_),
    .B(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__a221oi_1 _4971_ (.A1(_0383_),
    .A2(_0484_),
    .B1(_0622_),
    .B2(_0388_),
    .C1(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__and4_1 _4972_ (.A(_1662_),
    .B(_1666_),
    .C(_1669_),
    .D(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__o22ai_2 _4973_ (.A1(_0571_),
    .A2(_0450_),
    .B1(_0570_),
    .B2(_0454_),
    .Y(_1675_));
 sky130_fd_sc_hd__a221oi_2 _4974_ (.A1(_2904_),
    .A2(_0930_),
    .B1(_0447_),
    .B2(_0931_),
    .C1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__inv_2 _4975_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1677_));
 sky130_fd_sc_hd__o22ai_1 _4976_ (.A1(_1677_),
    .A2(_0464_),
    .B1(_1060_),
    .B2(_0467_),
    .Y(_1678_));
 sky130_fd_sc_hd__a221oi_1 _4977_ (.A1(_2962_),
    .A2(_0936_),
    .B1(_2817_),
    .B2(_0937_),
    .C1(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(_0438_),
    .B(_2865_),
    .Y(_1680_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_0442_),
    .B(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_1681_));
 sky130_fd_sc_hd__nand2_1 _4980_ (.A(_1680_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__a221oi_1 _4981_ (.A1(_2908_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_3083_),
    .C1(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__nand2_1 _4982_ (.A(_0420_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_1 _4983_ (.A(_0424_),
    .B(_0379_),
    .Y(_1685_));
 sky130_fd_sc_hd__nand2_1 _4984_ (.A(_1684_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__a221oi_1 _4985_ (.A1(_0414_),
    .A2(_0422_),
    .B1(_0417_),
    .B2(_3064_),
    .C1(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__and4_1 _4986_ (.A(_1676_),
    .B(_1679_),
    .C(_1683_),
    .D(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__and4_1 _4987_ (.A(_1648_),
    .B(_1659_),
    .C(_1674_),
    .D(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__nand3_2 _4988_ (.A(_1633_),
    .B(_3113_),
    .C(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__o21a_1 _4989_ (.A1(_0647_),
    .A2(_3112_),
    .B1(_2775_),
    .X(_1691_));
 sky130_fd_sc_hd__a22o_1 _4990_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B1(_1690_),
    .B2(_1691_),
    .X(_0288_));
 sky130_fd_sc_hd__a22o_1 _4991_ (.A1(_2853_),
    .A2(_2998_),
    .B1(_2856_),
    .B2(_0648_),
    .X(_1692_));
 sky130_fd_sc_hd__a221oi_1 _4992_ (.A1(_0566_),
    .A2(_0824_),
    .B1(_0507_),
    .B2(_0825_),
    .C1(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_1 _4993_ (.A(_2837_),
    .B(_0326_),
    .Y(_1694_));
 sky130_fd_sc_hd__nand2_1 _4994_ (.A(_2844_),
    .B(_2788_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_1694_),
    .B(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__a221oi_2 _4996_ (.A1(_2880_),
    .A2(_2826_),
    .B1(_2786_),
    .B2(_2831_),
    .C1(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__inv_2 _4997_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_1 _4998_ (.A(_2879_),
    .B(_2800_),
    .Y(_1699_));
 sky130_fd_sc_hd__o221a_1 _4999_ (.A1(_1098_),
    .A2(_2869_),
    .B1(_1698_),
    .B2(_2875_),
    .C1(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__nand2_1 _5000_ (.A(_2889_),
    .B(_2794_),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _5001_ (.A(_2893_),
    .B(_0589_),
    .Y(_1702_));
 sky130_fd_sc_hd__nand2_1 _5002_ (.A(_1701_),
    .B(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__a221oi_1 _5003_ (.A1(_2884_),
    .A2(_2790_),
    .B1(_2887_),
    .B2(_2812_),
    .C1(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__and4_1 _5004_ (.A(_1693_),
    .B(_1697_),
    .C(_1700_),
    .D(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__o22ai_1 _5005_ (.A1(_0932_),
    .A2(_2910_),
    .B1(_0570_),
    .B2(_2915_),
    .Y(_1706_));
 sky130_fd_sc_hd__a221oi_1 _5006_ (.A1(_3017_),
    .A2(_2902_),
    .B1(_0338_),
    .B2(_2906_),
    .C1(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__nand2_1 _5007_ (.A(_2924_),
    .B(_0524_),
    .Y(_1708_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_2927_),
    .B(_2810_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_1 _5009_ (.A(_1708_),
    .B(_1709_),
    .Y(_1710_));
 sky130_fd_sc_hd__a221oi_1 _5010_ (.A1(_2919_),
    .A2(_2777_),
    .B1(_2922_),
    .B2(_3078_),
    .C1(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__nand2_1 _5011_ (.A(_2943_),
    .B(_2808_),
    .Y(_1712_));
 sky130_fd_sc_hd__nand2_1 _5012_ (.A(_2947_),
    .B(_0436_),
    .Y(_1713_));
 sky130_fd_sc_hd__nand2_1 _5013_ (.A(_1712_),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__a221oi_1 _5014_ (.A1(_0471_),
    .A2(_2938_),
    .B1(_2940_),
    .B2(_2814_),
    .C1(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__nand2_1 _5015_ (.A(_2960_),
    .B(_0695_),
    .Y(_1716_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(_2964_),
    .B(_2792_),
    .Y(_1717_));
 sky130_fd_sc_hd__nand2_1 _5017_ (.A(_1716_),
    .B(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__a221oi_1 _5018_ (.A1(_3013_),
    .A2(_2954_),
    .B1(_0768_),
    .B2(_2958_),
    .C1(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__and4_1 _5019_ (.A(_1707_),
    .B(_1711_),
    .C(_1715_),
    .D(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__nand2_1 _5020_ (.A(_2985_),
    .B(_0384_),
    .Y(_1721_));
 sky130_fd_sc_hd__o21ai_1 _5021_ (.A1(_0741_),
    .A2(_2983_),
    .B1(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__a221oi_1 _5022_ (.A1(_2899_),
    .A2(_2975_),
    .B1(_3005_),
    .B2(_2980_),
    .C1(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__or2_1 _5023_ (.A(_3084_),
    .B(_0858_),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(_2996_),
    .B(_2977_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _5025_ (.A(_3000_),
    .B(_2846_),
    .Y(_1726_));
 sky130_fd_sc_hd__o2111a_1 _5026_ (.A1(_2909_),
    .A2(_2992_),
    .B1(_1724_),
    .C1(_1725_),
    .D1(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__o22ai_1 _5027_ (.A1(_1249_),
    .A2(_3015_),
    .B1(_0481_),
    .B2(_3021_),
    .Y(_1728_));
 sky130_fd_sc_hd__a221oi_1 _5028_ (.A1(_3050_),
    .A2(_3007_),
    .B1(_0358_),
    .B2(_3011_),
    .C1(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hd__nand2_1 _5029_ (.A(_3034_),
    .B(_2886_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_3038_),
    .B(_3098_),
    .Y(_1731_));
 sky130_fd_sc_hd__nand2_1 _5031_ (.A(_1730_),
    .B(_1731_),
    .Y(_1732_));
 sky130_fd_sc_hd__a221oi_1 _5032_ (.A1(_3027_),
    .A2(_0596_),
    .B1(_0410_),
    .B2(_3032_),
    .C1(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__and4_1 _5033_ (.A(_1723_),
    .B(_1727_),
    .C(_1729_),
    .D(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(_3051_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_3056_),
    .B(_0364_),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2_1 _5036_ (.A(_1735_),
    .B(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__a221oi_2 _5037_ (.A1(_3118_),
    .A2(_3046_),
    .B1(_3048_),
    .B2(_0510_),
    .C1(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__nand2_1 _5038_ (.A(_3068_),
    .B(_0591_),
    .Y(_1739_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(_3071_),
    .B(_0550_),
    .Y(_1740_));
 sky130_fd_sc_hd__nand2_1 _5040_ (.A(_1739_),
    .B(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hd__a221oi_1 _5041_ (.A1(_3062_),
    .A2(_0379_),
    .B1(_3065_),
    .B2(_0574_),
    .C1(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__nand2_1 _5042_ (.A(_3087_),
    .B(_2971_),
    .Y(_1743_));
 sky130_fd_sc_hd__o21ai_1 _5043_ (.A1(_0933_),
    .A2(_3085_),
    .B1(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__a221oi_1 _5044_ (.A1(_3076_),
    .A2(_3134_),
    .B1(_0323_),
    .B2(_3081_),
    .C1(_1744_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2_1 _5045_ (.A(_3099_),
    .B(_3104_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5046_ (.A(_3102_),
    .B(_0791_),
    .Y(_1747_));
 sky130_fd_sc_hd__nand2_1 _5047_ (.A(_1746_),
    .B(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__a221oi_1 _5048_ (.A1(_0513_),
    .A2(_3094_),
    .B1(_3096_),
    .B2(_3002_),
    .C1(_1748_),
    .Y(_1749_));
 sky130_fd_sc_hd__and4_1 _5049_ (.A(_1738_),
    .B(_1742_),
    .C(_1745_),
    .D(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__and4_1 _5050_ (.A(_1705_),
    .B(_1720_),
    .C(_1734_),
    .D(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__nand2_1 _5051_ (.A(_3126_),
    .B(_0395_),
    .Y(_1752_));
 sky130_fd_sc_hd__o21ai_1 _5052_ (.A1(_1645_),
    .A2(_3124_),
    .B1(_1752_),
    .Y(_1753_));
 sky130_fd_sc_hd__a221oi_1 _5053_ (.A1(_3079_),
    .A2(_3117_),
    .B1(_3067_),
    .B2(_3121_),
    .C1(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__or2_1 _5054_ (.A(_0656_),
    .B(_3136_),
    .X(_1755_));
 sky130_fd_sc_hd__or2_1 _5055_ (.A(_2913_),
    .B(_3140_),
    .X(_1756_));
 sky130_fd_sc_hd__nand2_1 _5056_ (.A(_3143_),
    .B(_0475_),
    .Y(_1757_));
 sky130_fd_sc_hd__o2111a_1 _5057_ (.A1(_1406_),
    .A2(_3132_),
    .B1(_1755_),
    .C1(_1756_),
    .D1(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__nand2_1 _5058_ (.A(_0324_),
    .B(_0595_),
    .Y(_1759_));
 sky130_fd_sc_hd__nand2_1 _5059_ (.A(_0328_),
    .B(_0451_),
    .Y(_1760_));
 sky130_fd_sc_hd__nand2_1 _5060_ (.A(_1759_),
    .B(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__a221oi_2 _5061_ (.A1(_3092_),
    .A2(_3149_),
    .B1(_3151_),
    .B2(_2932_),
    .C1(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__inv_2 _5062_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_1763_));
 sky130_fd_sc_hd__o22ai_1 _5063_ (.A1(_1763_),
    .A2(_0344_),
    .B1(_3122_),
    .B2(_0348_),
    .Y(_1764_));
 sky130_fd_sc_hd__a221oi_1 _5064_ (.A1(_0484_),
    .A2(_0336_),
    .B1(_0884_),
    .B2(_0340_),
    .C1(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__and4_1 _5065_ (.A(_1754_),
    .B(_1758_),
    .C(_1762_),
    .D(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__o22ai_1 _5066_ (.A1(_0676_),
    .A2(_0908_),
    .B1(_3131_),
    .B2(_0909_),
    .Y(_1767_));
 sky130_fd_sc_hd__a221oi_1 _5067_ (.A1(_3044_),
    .A2(_0906_),
    .B1(_3058_),
    .B2(_0907_),
    .C1(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__o22ai_1 _5068_ (.A1(_0816_),
    .A2(_0482_),
    .B1(_0606_),
    .B2(_0486_),
    .Y(_1769_));
 sky130_fd_sc_hd__a221oi_1 _5069_ (.A1(_0622_),
    .A2(_0477_),
    .B1(_0352_),
    .B2(_2757_),
    .C1(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__o22ai_1 _5070_ (.A1(_1219_),
    .A2(_0503_),
    .B1(_1677_),
    .B2(_0915_),
    .Y(_1771_));
 sky130_fd_sc_hd__a22o_1 _5071_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .B1(_0918_),
    .B2(_2802_),
    .X(_1772_));
 sky130_fd_sc_hd__nor2_1 _5072_ (.A(_1771_),
    .B(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__o22ai_1 _5073_ (.A1(_0342_),
    .A2(_0922_),
    .B1(_1043_),
    .B2(_0923_),
    .Y(_1774_));
 sky130_fd_sc_hd__a22o_1 _5074_ (.A1(_0925_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .B1(_0926_),
    .B2(_0647_),
    .X(_1775_));
 sky130_fd_sc_hd__nor2_1 _5075_ (.A(_1774_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__and4_1 _5076_ (.A(_1768_),
    .B(_1770_),
    .C(_1773_),
    .D(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__nand2_1 _5077_ (.A(_0372_),
    .B(_0439_),
    .Y(_1778_));
 sky130_fd_sc_hd__o21ai_1 _5078_ (.A1(_0801_),
    .A2(_0369_),
    .B1(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__a221oi_2 _5079_ (.A1(_2962_),
    .A2(_0378_),
    .B1(_0649_),
    .B2(_0375_),
    .C1(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__nand2_1 _5080_ (.A(_0359_),
    .B(_0416_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_1 _5081_ (.A(_0362_),
    .B(_0584_),
    .Y(_1782_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_1781_),
    .B(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__a221oi_2 _5083_ (.A1(_0707_),
    .A2(_0354_),
    .B1(_0356_),
    .B2(_3053_),
    .C1(_1783_),
    .Y(_1784_));
 sky130_fd_sc_hd__a22o_1 _5084_ (.A1(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_1785_));
 sky130_fd_sc_hd__a22o_1 _5085_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .B1(_0409_),
    .B2(_0651_),
    .X(_1786_));
 sky130_fd_sc_hd__nor2_1 _5086_ (.A(_1785_),
    .B(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__nand2_1 _5087_ (.A(_0390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1788_));
 sky130_fd_sc_hd__nand2_1 _5088_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_1789_));
 sky130_fd_sc_hd__nand2_1 _5089_ (.A(_1788_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__a221oi_1 _5090_ (.A1(_0383_),
    .A2(_0345_),
    .B1(_3029_),
    .B2(_0388_),
    .C1(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__and4_1 _5091_ (.A(_1780_),
    .B(_1784_),
    .C(_1787_),
    .D(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__o22ai_1 _5092_ (.A1(_0725_),
    .A2(_0449_),
    .B1(_0724_),
    .B2(_0453_),
    .Y(_1793_));
 sky130_fd_sc_hd__a221oi_2 _5093_ (.A1(_0447_),
    .A2(_0930_),
    .B1(_2987_),
    .B2(_0931_),
    .C1(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__o22ai_1 _5094_ (.A1(_2868_),
    .A2(_0463_),
    .B1(_1181_),
    .B2(_0466_),
    .Y(_1795_));
 sky130_fd_sc_hd__a221oi_1 _5095_ (.A1(_2817_),
    .A2(_0936_),
    .B1(_2865_),
    .B2(_0937_),
    .C1(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__nand2_1 _5096_ (.A(_0437_),
    .B(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_1797_));
 sky130_fd_sc_hd__nand2_1 _5097_ (.A(_0441_),
    .B(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1798_));
 sky130_fd_sc_hd__nand2_1 _5098_ (.A(_1797_),
    .B(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__a221oi_1 _5099_ (.A1(_2952_),
    .A2(_0432_),
    .B1(_0434_),
    .B2(_0457_),
    .C1(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__nand2_1 _5100_ (.A(_0420_),
    .B(_0746_),
    .Y(_1801_));
 sky130_fd_sc_hd__nand2_1 _5101_ (.A(_0424_),
    .B(_0631_),
    .Y(_1802_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(_1801_),
    .B(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__a221oi_1 _5103_ (.A1(_0414_),
    .A2(_3030_),
    .B1(_0417_),
    .B2(_0426_),
    .C1(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__and4_1 _5104_ (.A(_1794_),
    .B(_1796_),
    .C(_1800_),
    .D(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__and4_1 _5105_ (.A(_1766_),
    .B(_1777_),
    .C(_1792_),
    .D(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__nand3_1 _5106_ (.A(_1751_),
    .B(_0525_),
    .C(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__o21a_1 _5107_ (.A1(_0330_),
    .A2(_3112_),
    .B1(_2775_),
    .X(_1808_));
 sky130_fd_sc_hd__a22o_1 _5108_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .B1(_1807_),
    .B2(_1808_),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_1 _5109_ (.A1(_2853_),
    .A2(_0566_),
    .B1(_2856_),
    .B2(_2998_),
    .X(_1809_));
 sky130_fd_sc_hd__a221oi_1 _5110_ (.A1(_2777_),
    .A2(_0825_),
    .B1(_0430_),
    .B2(_0824_),
    .C1(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__nand2_1 _5111_ (.A(_2837_),
    .B(_3017_),
    .Y(_1811_));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(_2844_),
    .B(_2790_),
    .Y(_1812_));
 sky130_fd_sc_hd__nand2_1 _5113_ (.A(_1811_),
    .B(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__a221oi_2 _5114_ (.A1(_0507_),
    .A2(_2826_),
    .B1(_2788_),
    .B2(_2831_),
    .C1(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_2878_),
    .B(_2802_),
    .Y(_1815_));
 sky130_fd_sc_hd__o21ai_1 _5116_ (.A1(_1219_),
    .A2(_2870_),
    .B1(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__a31oi_1 _5117_ (.A1(_2808_),
    .A2(_2860_),
    .A3(_2874_),
    .B1(_1816_),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _5118_ (.A(_2889_),
    .B(_2796_),
    .Y(_1818_));
 sky130_fd_sc_hd__nand2_1 _5119_ (.A(_2893_),
    .B(_0591_),
    .Y(_1819_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_1818_),
    .B(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__a221oi_1 _5121_ (.A1(_2884_),
    .A2(_2792_),
    .B1(_2887_),
    .B2(_2814_),
    .C1(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__and4_1 _5122_ (.A(_1810_),
    .B(_1814_),
    .C(_1817_),
    .D(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__o22ai_1 _5123_ (.A1(_3014_),
    .A2(_2910_),
    .B1(_0724_),
    .B2(_2915_),
    .Y(_1823_));
 sky130_fd_sc_hd__a221oi_1 _5124_ (.A1(_0338_),
    .A2(_2902_),
    .B1(_0334_),
    .B2(_2906_),
    .C1(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__nand2_1 _5125_ (.A(_2924_),
    .B(_3078_),
    .Y(_1825_));
 sky130_fd_sc_hd__nand2_1 _5126_ (.A(_2927_),
    .B(_2812_),
    .Y(_1826_));
 sky130_fd_sc_hd__nand2_1 _5127_ (.A(_1825_),
    .B(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__a221oi_1 _5128_ (.A1(_2919_),
    .A2(_2786_),
    .B1(_2922_),
    .B2(_0589_),
    .C1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand2_1 _5129_ (.A(_2943_),
    .B(_2810_),
    .Y(_1829_));
 sky130_fd_sc_hd__nand2_1 _5130_ (.A(_2947_),
    .B(_0648_),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _5131_ (.A(_1829_),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__a221oi_1 _5132_ (.A1(_0439_),
    .A2(_2938_),
    .B1(_2940_),
    .B2(_0524_),
    .C1(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(_2960_),
    .B(_2880_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _5134_ (.A(_2964_),
    .B(_2794_),
    .Y(_1834_));
 sky130_fd_sc_hd__nand2_1 _5135_ (.A(_1833_),
    .B(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__a221oi_1 _5136_ (.A1(_2956_),
    .A2(_2954_),
    .B1(_3092_),
    .B2(_2958_),
    .C1(_1835_),
    .Y(_1836_));
 sky130_fd_sc_hd__and4_1 _5137_ (.A(_1824_),
    .B(_1828_),
    .C(_1832_),
    .D(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__nand2_1 _5138_ (.A(_2985_),
    .B(_3050_),
    .Y(_1838_));
 sky130_fd_sc_hd__o21ai_1 _5139_ (.A1(_0880_),
    .A2(_2983_),
    .B1(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__a221oi_1 _5140_ (.A1(_2904_),
    .A2(_2975_),
    .B1(_3009_),
    .B2(_2980_),
    .C1(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__or2_1 _5141_ (.A(_0590_),
    .B(_0858_),
    .X(_1841_));
 sky130_fd_sc_hd__nand2_1 _5142_ (.A(_2996_),
    .B(_2908_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _5143_ (.A(_3000_),
    .B(_2886_),
    .Y(_1843_));
 sky130_fd_sc_hd__o2111a_1 _5144_ (.A1(_0543_),
    .A2(_2992_),
    .B1(_1841_),
    .C1(_1842_),
    .D1(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__o22ai_1 _5145_ (.A1(_1370_),
    .A2(_3015_),
    .B1(_0492_),
    .B2(_3021_),
    .Y(_1845_));
 sky130_fd_sc_hd__a221oi_1 _5146_ (.A1(_0358_),
    .A2(_3007_),
    .B1(_0623_),
    .B2(_3011_),
    .C1(_1845_),
    .Y(_1846_));
 sky130_fd_sc_hd__nand2_1 _5147_ (.A(_3034_),
    .B(_2966_),
    .Y(_1847_));
 sky130_fd_sc_hd__nand2_1 _5148_ (.A(_3038_),
    .B(_0596_),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_1847_),
    .B(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__a221oi_1 _5150_ (.A1(_3027_),
    .A2(_0746_),
    .B1(_3104_),
    .B2(_3032_),
    .C1(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__and4_1 _5151_ (.A(_1840_),
    .B(_1844_),
    .C(_1846_),
    .D(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__nand2_1 _5152_ (.A(_3051_),
    .B(_3118_),
    .Y(_1852_));
 sky130_fd_sc_hd__nand2_1 _5153_ (.A(_3056_),
    .B(_0391_),
    .Y(_1853_));
 sky130_fd_sc_hd__nand2_1 _5154_ (.A(_1852_),
    .B(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__a221oi_2 _5155_ (.A1(_0364_),
    .A2(_3046_),
    .B1(_3048_),
    .B2(_3053_),
    .C1(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__nand2_1 _5156_ (.A(_3068_),
    .B(_0436_),
    .Y(_1856_));
 sky130_fd_sc_hd__nand2_1 _5157_ (.A(_3071_),
    .B(_0707_),
    .Y(_1857_));
 sky130_fd_sc_hd__nand2_1 _5158_ (.A(_1856_),
    .B(_1857_),
    .Y(_1858_));
 sky130_fd_sc_hd__a221oi_1 _5159_ (.A1(_3062_),
    .A2(_0631_),
    .B1(_3065_),
    .B2(_3064_),
    .C1(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__nand2_1 _5160_ (.A(_3087_),
    .B(_3083_),
    .Y(_1860_));
 sky130_fd_sc_hd__o21ai_1 _5161_ (.A1(_0448_),
    .A2(_3085_),
    .B1(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hd__a221oi_2 _5162_ (.A1(_3076_),
    .A2(_2971_),
    .B1(_0613_),
    .B2(_3081_),
    .C1(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__nand2_1 _5163_ (.A(_3099_),
    .B(_0379_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand2_1 _5164_ (.A(_3102_),
    .B(_2962_),
    .Y(_1864_));
 sky130_fd_sc_hd__nand2_1 _5165_ (.A(_1863_),
    .B(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__a221oi_1 _5166_ (.A1(_3114_),
    .A2(_3094_),
    .B1(_3096_),
    .B2(_3036_),
    .C1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__and4_1 _5167_ (.A(_1855_),
    .B(_1859_),
    .C(_1862_),
    .D(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__and4_1 _5168_ (.A(_1822_),
    .B(_1837_),
    .C(_1851_),
    .D(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__nand2_1 _5169_ (.A(_3125_),
    .B(_0479_),
    .Y(_1869_));
 sky130_fd_sc_hd__o21ai_1 _5170_ (.A1(_1763_),
    .A2(_3123_),
    .B1(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__a221oi_1 _5171_ (.A1(_0395_),
    .A2(_3116_),
    .B1(_0584_),
    .B2(_3120_),
    .C1(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__or2_1 _5172_ (.A(_0796_),
    .B(_3136_),
    .X(_1872_));
 sky130_fd_sc_hd__or2_1 _5173_ (.A(_0452_),
    .B(_3140_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2_1 _5174_ (.A(_3143_),
    .B(_0385_),
    .Y(_1874_));
 sky130_fd_sc_hd__o2111a_1 _5175_ (.A1(_1527_),
    .A2(_3132_),
    .B1(_1872_),
    .C1(_1873_),
    .D1(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__nand2_1 _5176_ (.A(_0324_),
    .B(_0745_),
    .Y(_1876_));
 sky130_fd_sc_hd__nand2_1 _5177_ (.A(_0328_),
    .B(_2839_),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(_1876_),
    .B(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__a221oi_2 _5179_ (.A1(_0595_),
    .A2(_3149_),
    .B1(_3151_),
    .B2(_0550_),
    .C1(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__inv_2 _5180_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_1880_));
 sky130_fd_sc_hd__o22ai_1 _5181_ (.A1(_1880_),
    .A2(_0343_),
    .B1(_0342_),
    .B2(_0347_),
    .Y(_1881_));
 sky130_fd_sc_hd__a221oi_1 _5182_ (.A1(_0345_),
    .A2(_0336_),
    .B1(_0484_),
    .B2(_0340_),
    .C1(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__and4_1 _5183_ (.A(_1871_),
    .B(_1875_),
    .C(_1879_),
    .D(_1882_),
    .X(_1883_));
 sky130_fd_sc_hd__o22ai_1 _5184_ (.A1(_0816_),
    .A2(_0908_),
    .B1(_0606_),
    .B2(_0909_),
    .Y(_1884_));
 sky130_fd_sc_hd__a221oi_1 _5185_ (.A1(_3058_),
    .A2(_0906_),
    .B1(_0513_),
    .B2(_0907_),
    .C1(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__o22ai_1 _5186_ (.A1(_3131_),
    .A2(_0482_),
    .B1(_3122_),
    .B2(_0486_),
    .Y(_1886_));
 sky130_fd_sc_hd__a221oi_1 _5187_ (.A1(_3029_),
    .A2(_0477_),
    .B1(_0622_),
    .B2(_2757_),
    .C1(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__o22ai_1 _5188_ (.A1(_1340_),
    .A2(_0503_),
    .B1(_2868_),
    .B2(_0915_),
    .Y(_1888_));
 sky130_fd_sc_hd__a22o_1 _5189_ (.A1(_0917_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .B1(_0918_),
    .B2(_2804_),
    .X(_1889_));
 sky130_fd_sc_hd__nor2_1 _5190_ (.A(_1888_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__o22ai_2 _5191_ (.A1(_0618_),
    .A2(_0922_),
    .B1(_1164_),
    .B2(_0923_),
    .Y(_1891_));
 sky130_fd_sc_hd__a22o_1 _5192_ (.A1(_0925_),
    .A2(_0647_),
    .B1(_0926_),
    .B2(_0330_),
    .X(_1892_));
 sky130_fd_sc_hd__nor2_1 _5193_ (.A(_1891_),
    .B(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__and4_1 _5194_ (.A(_1885_),
    .B(_1887_),
    .C(_1890_),
    .D(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__nand2_1 _5195_ (.A(_0372_),
    .B(_0649_),
    .Y(_1895_));
 sky130_fd_sc_hd__o21ai_1 _5196_ (.A1(_0939_),
    .A2(_0369_),
    .B1(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__a221oi_2 _5197_ (.A1(_2817_),
    .A2(_0378_),
    .B1(_3002_),
    .B2(_0375_),
    .C1(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__nand2_1 _5198_ (.A(_0359_),
    .B(_3067_),
    .Y(_1898_));
 sky130_fd_sc_hd__nand2_1 _5199_ (.A(_0362_),
    .B(_0419_),
    .Y(_1899_));
 sky130_fd_sc_hd__nand2_1 _5200_ (.A(_1898_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__a221oi_2 _5201_ (.A1(_3098_),
    .A2(_0354_),
    .B1(_0356_),
    .B2(_3044_),
    .C1(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__a22o_1 _5202_ (.A1(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .A2(_0401_),
    .B1(_0404_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_1902_));
 sky130_fd_sc_hd__a22o_1 _5203_ (.A1(_0407_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .B1(_0409_),
    .B2(_0791_),
    .X(_1903_));
 sky130_fd_sc_hd__nor2_1 _5204_ (.A(_1902_),
    .B(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__nand2_1 _5205_ (.A(_0390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_0394_),
    .B(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _5207_ (.A(_1905_),
    .B(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__a221oi_1 _5208_ (.A1(_0383_),
    .A2(_0510_),
    .B1(_0422_),
    .B2(_0388_),
    .C1(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__and4_1 _5209_ (.A(_1897_),
    .B(_1901_),
    .C(_1904_),
    .D(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__o22ai_2 _5210_ (.A1(_0864_),
    .A2(_0449_),
    .B1(_0863_),
    .B2(_0453_),
    .Y(_1910_));
 sky130_fd_sc_hd__a221oi_2 _5211_ (.A1(_2987_),
    .A2(_0930_),
    .B1(_3005_),
    .B2(_0931_),
    .C1(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__o22ai_1 _5212_ (.A1(_0501_),
    .A2(_0463_),
    .B1(_1302_),
    .B2(_0466_),
    .Y(_1912_));
 sky130_fd_sc_hd__a221oi_1 _5213_ (.A1(_2865_),
    .A2(_0936_),
    .B1(_2921_),
    .B2(_0937_),
    .C1(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__nand2_1 _5214_ (.A(_0437_),
    .B(_2828_),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _5215_ (.A(_0441_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1915_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_1914_),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__a221oi_1 _5217_ (.A1(_2912_),
    .A2(_0432_),
    .B1(_0434_),
    .B2(_0459_),
    .C1(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(_0420_),
    .B(_0410_),
    .Y(_1918_));
 sky130_fd_sc_hd__nand2_1 _5219_ (.A(_0424_),
    .B(_0471_),
    .Y(_1919_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(_1918_),
    .B(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__a221oi_1 _5221_ (.A1(_0414_),
    .A2(_0574_),
    .B1(_0417_),
    .B2(_2932_),
    .C1(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__and4_1 _5222_ (.A(_1911_),
    .B(_1913_),
    .C(_1917_),
    .D(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__and4_1 _5223_ (.A(_1883_),
    .B(_1894_),
    .C(_1909_),
    .D(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__nand3_1 _5224_ (.A(_1868_),
    .B(_0525_),
    .C(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__o21a_1 _5225_ (.A1(_3134_),
    .A2(_3112_),
    .B1(_2775_),
    .X(_1925_));
 sky130_fd_sc_hd__a22o_1 _5226_ (.A1(_2816_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .B1(_1924_),
    .B2(_1925_),
    .X(_0286_));
 sky130_fd_sc_hd__inv_2 _5227_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_1926_));
 sky130_fd_sc_hd__a22o_1 _5228_ (.A1(_0574_),
    .A2(_0401_),
    .B1(_0404_),
    .B2(_2932_),
    .X(_1927_));
 sky130_fd_sc_hd__a221oi_1 _5229_ (.A1(_0791_),
    .A2(_0407_),
    .B1(_2962_),
    .B2(_0409_),
    .C1(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__nand2_1 _5230_ (.A(_0372_),
    .B(_3002_),
    .Y(_1929_));
 sky130_fd_sc_hd__o21ai_1 _5231_ (.A1(_0499_),
    .A2(_0369_),
    .B1(_1929_),
    .Y(_1930_));
 sky130_fd_sc_hd__a221oi_2 _5232_ (.A1(_2865_),
    .A2(_0378_),
    .B1(_3036_),
    .B2(_0375_),
    .C1(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_0390_),
    .B(_0613_),
    .Y(_1932_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(_0394_),
    .B(_0622_),
    .Y(_1933_));
 sky130_fd_sc_hd__nand2_1 _5235_ (.A(_1932_),
    .B(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__a221oi_1 _5236_ (.A1(_0383_),
    .A2(_3053_),
    .B1(_3030_),
    .B2(_0388_),
    .C1(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__nand2_1 _5237_ (.A(_0360_),
    .B(_0584_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _5238_ (.A(_0363_),
    .B(_0323_),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(_1936_),
    .B(_1937_),
    .Y(_1938_));
 sky130_fd_sc_hd__a221oi_1 _5240_ (.A1(_0596_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_3058_),
    .C1(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__and4_1 _5241_ (.A(_1928_),
    .B(_1931_),
    .C(_1935_),
    .D(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_3126_),
    .B(_0475_),
    .Y(_1941_));
 sky130_fd_sc_hd__o21ai_1 _5243_ (.A1(_1880_),
    .A2(_3124_),
    .B1(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__a221oi_1 _5244_ (.A1(_0479_),
    .A2(_3117_),
    .B1(_0419_),
    .B2(_3121_),
    .C1(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__or2_1 _5245_ (.A(_0933_),
    .B(_3137_),
    .X(_1944_));
 sky130_fd_sc_hd__or2_1 _5246_ (.A(_0656_),
    .B(_3141_),
    .X(_1945_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(_3144_),
    .B(_0634_),
    .Y(_1946_));
 sky130_fd_sc_hd__o2111a_1 _5248_ (.A1(_1645_),
    .A2(_3133_),
    .B1(_1944_),
    .C1(_1945_),
    .D1(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__nand2_1 _5249_ (.A(_0325_),
    .B(_0884_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand2_1 _5250_ (.A(_0329_),
    .B(_2899_),
    .Y(_1949_));
 sky130_fd_sc_hd__nand2_1 _5251_ (.A(_1948_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__a221oi_2 _5252_ (.A1(_0745_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0707_),
    .C1(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hd__inv_2 _5253_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1952_));
 sky130_fd_sc_hd__o22ai_1 _5254_ (.A1(_1952_),
    .A2(_0344_),
    .B1(_0618_),
    .B2(_0348_),
    .Y(_1953_));
 sky130_fd_sc_hd__a221oi_1 _5255_ (.A1(_0510_),
    .A2(_0337_),
    .B1(_0345_),
    .B2(_0341_),
    .C1(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__and4_1 _5256_ (.A(_1943_),
    .B(_1947_),
    .C(_1951_),
    .D(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__o22ai_1 _5257_ (.A1(_1007_),
    .A2(_0450_),
    .B1(_3018_),
    .B2(_0454_),
    .Y(_1956_));
 sky130_fd_sc_hd__a221oi_1 _5258_ (.A1(_3005_),
    .A2(_0930_),
    .B1(_3009_),
    .B2(_0931_),
    .C1(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__o22ai_1 _5259_ (.A1(_0671_),
    .A2(_0464_),
    .B1(_1423_),
    .B2(_0467_),
    .Y(_1958_));
 sky130_fd_sc_hd__a221oi_1 _5260_ (.A1(_2921_),
    .A2(_0936_),
    .B1(_2828_),
    .B2(_0937_),
    .C1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nand2_1 _5261_ (.A(_0438_),
    .B(_2846_),
    .Y(_1960_));
 sky130_fd_sc_hd__nand2_1 _5262_ (.A(_0442_),
    .B(_0537_),
    .Y(_1961_));
 sky130_fd_sc_hd__nand2_1 _5263_ (.A(_1960_),
    .B(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__a221oi_1 _5264_ (.A1(_0451_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_2977_),
    .C1(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_0421_),
    .B(_3104_),
    .Y(_1964_));
 sky130_fd_sc_hd__nand2_1 _5266_ (.A(_0425_),
    .B(_0439_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand2_1 _5267_ (.A(_1964_),
    .B(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__a221oi_1 _5268_ (.A1(_0415_),
    .A2(_3064_),
    .B1(_0418_),
    .B2(_0550_),
    .C1(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__and4_1 _5269_ (.A(_1957_),
    .B(_1959_),
    .C(_1963_),
    .D(_1967_),
    .X(_1968_));
 sky130_fd_sc_hd__o22ai_1 _5270_ (.A1(_3131_),
    .A2(_0908_),
    .B1(_3122_),
    .B2(_0909_),
    .Y(_1969_));
 sky130_fd_sc_hd__a221oi_1 _5271_ (.A1(_0513_),
    .A2(_0906_),
    .B1(_3114_),
    .B2(_0907_),
    .C1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__o22ai_2 _5272_ (.A1(_1461_),
    .A2(_0503_),
    .B1(_0501_),
    .B2(_0915_),
    .Y(_1971_));
 sky130_fd_sc_hd__a221oi_4 _5273_ (.A1(_2806_),
    .A2(_0918_),
    .B1(_2808_),
    .B2(_0917_),
    .C1(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__o22ai_1 _5274_ (.A1(_0606_),
    .A2(_0483_),
    .B1(_0342_),
    .B2(_0487_),
    .Y(_1973_));
 sky130_fd_sc_hd__a221oi_1 _5275_ (.A1(_0422_),
    .A2(_0478_),
    .B1(_3029_),
    .B2(_0480_),
    .C1(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__o22ai_1 _5276_ (.A1(_0764_),
    .A2(_0922_),
    .B1(_1285_),
    .B2(_0923_),
    .Y(_1975_));
 sky130_fd_sc_hd__a221oi_1 _5277_ (.A1(_0330_),
    .A2(_0925_),
    .B1(_3134_),
    .B2(_0926_),
    .C1(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__and4_1 _5278_ (.A(_1970_),
    .B(_1972_),
    .C(_1974_),
    .D(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__and4_1 _5279_ (.A(_1940_),
    .B(_1955_),
    .C(_1968_),
    .D(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__a22o_1 _5280_ (.A1(_2854_),
    .A2(_0430_),
    .B1(_2857_),
    .B2(_0566_),
    .X(_1979_));
 sky130_fd_sc_hd__a221oi_1 _5281_ (.A1(_2786_),
    .A2(_0825_),
    .B1(_0647_),
    .B2(_0824_),
    .C1(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _5282_ (.A(_2838_),
    .B(_0338_),
    .Y(_1981_));
 sky130_fd_sc_hd__nand2_1 _5283_ (.A(_2845_),
    .B(_2792_),
    .Y(_1982_));
 sky130_fd_sc_hd__nand2_1 _5284_ (.A(_1981_),
    .B(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__a221oi_1 _5285_ (.A1(_2777_),
    .A2(_2827_),
    .B1(_2790_),
    .B2(_2832_),
    .C1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__nand2_1 _5286_ (.A(_2879_),
    .B(_2804_),
    .Y(_1985_));
 sky130_fd_sc_hd__o21ai_1 _5287_ (.A1(_1340_),
    .A2(_2870_),
    .B1(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__a31oi_1 _5288_ (.A1(_2810_),
    .A2(_2860_),
    .A3(_2874_),
    .B1(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _5289_ (.A(_2890_),
    .B(_2798_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5290_ (.A(_2894_),
    .B(_0436_),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _5291_ (.A(_1988_),
    .B(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__a221oi_1 _5292_ (.A1(_2885_),
    .A2(_2794_),
    .B1(_2888_),
    .B2(_0524_),
    .C1(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__and4_1 _5293_ (.A(_1980_),
    .B(_1984_),
    .C(_1987_),
    .D(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__o22ai_1 _5294_ (.A1(_0570_),
    .A2(_2911_),
    .B1(_0863_),
    .B2(_2916_),
    .Y(_1993_));
 sky130_fd_sc_hd__a221oi_1 _5295_ (.A1(_0334_),
    .A2(_2903_),
    .B1(_0384_),
    .B2(_2907_),
    .C1(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__nand2_1 _5296_ (.A(_2925_),
    .B(_0589_),
    .Y(_1995_));
 sky130_fd_sc_hd__nand2_1 _5297_ (.A(_2928_),
    .B(_2814_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_1 _5298_ (.A(_1995_),
    .B(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__a221oi_1 _5299_ (.A1(_2920_),
    .A2(_2788_),
    .B1(_2923_),
    .B2(_0591_),
    .C1(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(_2944_),
    .B(_2812_),
    .Y(_1999_));
 sky130_fd_sc_hd__nand2_1 _5301_ (.A(_2948_),
    .B(_2998_),
    .Y(_2000_));
 sky130_fd_sc_hd__nand2_1 _5302_ (.A(_1999_),
    .B(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hd__a221oi_1 _5303_ (.A1(_0649_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_3078_),
    .C1(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__nand2_1 _5304_ (.A(_2961_),
    .B(_0507_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _5305_ (.A(_2965_),
    .B(_2796_),
    .Y(_2004_));
 sky130_fd_sc_hd__nand2_1 _5306_ (.A(_2003_),
    .B(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__a221oi_1 _5307_ (.A1(_3147_),
    .A2(_2955_),
    .B1(_0595_),
    .B2(_2959_),
    .C1(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__and4_1 _5308_ (.A(_1994_),
    .B(_1998_),
    .C(_2002_),
    .D(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__nand2_1 _5309_ (.A(_2986_),
    .B(_0358_),
    .Y(_2008_));
 sky130_fd_sc_hd__o21ai_1 _5310_ (.A1(_2909_),
    .A2(_2984_),
    .B1(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__a221oi_1 _5311_ (.A1(_0447_),
    .A2(_2976_),
    .B1(_3013_),
    .B2(_2981_),
    .C1(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__or2_1 _5312_ (.A(_0741_),
    .B(_0858_),
    .X(_2011_));
 sky130_fd_sc_hd__nand2_1 _5313_ (.A(_2997_),
    .B(_2952_),
    .Y(_2012_));
 sky130_fd_sc_hd__nand2_1 _5314_ (.A(_3001_),
    .B(_2966_),
    .Y(_2013_));
 sky130_fd_sc_hd__o2111a_1 _5315_ (.A1(_2913_),
    .A2(_2993_),
    .B1(_2011_),
    .C1(_2012_),
    .D1(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__o22ai_1 _5316_ (.A1(_1491_),
    .A2(_3016_),
    .B1(_0485_),
    .B2(_3022_),
    .Y(_2015_));
 sky130_fd_sc_hd__a221oi_2 _5317_ (.A1(_0623_),
    .A2(_3008_),
    .B1(_0768_),
    .B2(_3012_),
    .C1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _5318_ (.A(_3035_),
    .B(_2891_),
    .Y(_2017_));
 sky130_fd_sc_hd__nand2_1 _5319_ (.A(_3039_),
    .B(_0746_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand2_1 _5320_ (.A(_2017_),
    .B(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__a221oi_1 _5321_ (.A1(_3028_),
    .A2(_0410_),
    .B1(_0379_),
    .B2(_3033_),
    .C1(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__and4_1 _5322_ (.A(_2010_),
    .B(_2014_),
    .C(_2016_),
    .D(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__nand2_1 _5323_ (.A(_3052_),
    .B(_0364_),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_1 _5324_ (.A(_3057_),
    .B(_3079_),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(_2022_),
    .B(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__a221oi_1 _5326_ (.A1(_0391_),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_3044_),
    .C1(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _5327_ (.A(_3069_),
    .B(_0648_),
    .Y(_2026_));
 sky130_fd_sc_hd__nand2_1 _5328_ (.A(_3072_),
    .B(_3098_),
    .Y(_2027_));
 sky130_fd_sc_hd__nand2_1 _5329_ (.A(_2026_),
    .B(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__a221oi_1 _5330_ (.A1(_3063_),
    .A2(_0471_),
    .B1(_3066_),
    .B2(_0426_),
    .C1(_2028_),
    .Y(_2029_));
 sky130_fd_sc_hd__nand2_1 _5331_ (.A(_3088_),
    .B(_0457_),
    .Y(_2030_));
 sky130_fd_sc_hd__o21ai_1 _5332_ (.A1(_0655_),
    .A2(_3086_),
    .B1(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__a221oi_1 _5333_ (.A1(_3077_),
    .A2(_3083_),
    .B1(_0352_),
    .B2(_3082_),
    .C1(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__nand2_1 _5334_ (.A(_3100_),
    .B(_0631_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand2_1 _5335_ (.A(_3103_),
    .B(_2817_),
    .Y(_2034_));
 sky130_fd_sc_hd__nand2_1 _5336_ (.A(_2033_),
    .B(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__a221oi_1 _5337_ (.A1(_3127_),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0443_),
    .C1(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__and4_1 _5338_ (.A(_2025_),
    .B(_2029_),
    .C(_2032_),
    .D(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__and4_1 _5339_ (.A(_1992_),
    .B(_2007_),
    .C(_2021_),
    .D(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__nand3_2 _5340_ (.A(_1978_),
    .B(_2038_),
    .C(_3113_),
    .Y(_2039_));
 sky130_fd_sc_hd__o21a_1 _5341_ (.A1(_2971_),
    .A2(_0525_),
    .B1(_2776_),
    .X(_2040_));
 sky130_fd_sc_hd__nand2_1 _5342_ (.A(_2039_),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__o21ai_1 _5343_ (.A1(_2776_),
    .A2(_1926_),
    .B1(_2041_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _5344_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2042_));
 sky130_fd_sc_hd__a22o_1 _5345_ (.A1(_3064_),
    .A2(_0401_),
    .B1(_0404_),
    .B2(_0550_),
    .X(_2043_));
 sky130_fd_sc_hd__a221oi_1 _5346_ (.A1(_2962_),
    .A2(_0407_),
    .B1(_2817_),
    .B2(_0409_),
    .C1(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__nand2_1 _5347_ (.A(_0372_),
    .B(_3036_),
    .Y(_2045_));
 sky130_fd_sc_hd__o21ai_1 _5348_ (.A1(_0462_),
    .A2(_0369_),
    .B1(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__a221oi_2 _5349_ (.A1(_0443_),
    .A2(_0375_),
    .B1(_2921_),
    .B2(_0378_),
    .C1(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__nand2_1 _5350_ (.A(_0390_),
    .B(_0352_),
    .Y(_2048_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(_0394_),
    .B(_3029_),
    .Y(_2049_));
 sky130_fd_sc_hd__nand2_1 _5352_ (.A(_2048_),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__a221oi_1 _5353_ (.A1(_0383_),
    .A2(_3044_),
    .B1(_0574_),
    .B2(_0388_),
    .C1(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__nand2_1 _5354_ (.A(_0360_),
    .B(_0419_),
    .Y(_2052_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_0363_),
    .B(_0613_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _5356_ (.A(_2052_),
    .B(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__a221oi_1 _5357_ (.A1(_0746_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_0513_),
    .C1(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__and4_1 _5358_ (.A(_2044_),
    .B(_2047_),
    .C(_2051_),
    .D(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__nand2_1 _5359_ (.A(_3126_),
    .B(_0385_),
    .Y(_2057_));
 sky130_fd_sc_hd__o21ai_1 _5360_ (.A1(_1952_),
    .A2(_3124_),
    .B1(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__a221oi_1 _5361_ (.A1(_0475_),
    .A2(_3117_),
    .B1(_0323_),
    .B2(_3121_),
    .C1(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__or2_1 _5362_ (.A(_0448_),
    .B(_3137_),
    .X(_2060_));
 sky130_fd_sc_hd__or2_1 _5363_ (.A(_0796_),
    .B(_3141_),
    .X(_2061_));
 sky130_fd_sc_hd__nand2_1 _5364_ (.A(_3144_),
    .B(_0416_),
    .Y(_2062_));
 sky130_fd_sc_hd__o2111a_1 _5365_ (.A1(_1763_),
    .A2(_3133_),
    .B1(_2060_),
    .C1(_2061_),
    .D1(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__nand2_1 _5366_ (.A(_0325_),
    .B(_0484_),
    .Y(_2064_));
 sky130_fd_sc_hd__nand2_1 _5367_ (.A(_0329_),
    .B(_2904_),
    .Y(_2065_));
 sky130_fd_sc_hd__nand2_1 _5368_ (.A(_2064_),
    .B(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__a221oi_2 _5369_ (.A1(_0884_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_3098_),
    .C1(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__inv_2 _5370_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_2068_));
 sky130_fd_sc_hd__o22ai_1 _5371_ (.A1(_2068_),
    .A2(_0344_),
    .B1(_0764_),
    .B2(_0348_),
    .Y(_2069_));
 sky130_fd_sc_hd__a221oi_1 _5372_ (.A1(_3053_),
    .A2(_0337_),
    .B1(_0510_),
    .B2(_0341_),
    .C1(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__and4_1 _5373_ (.A(_2059_),
    .B(_2063_),
    .C(_2067_),
    .D(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__o22ai_1 _5374_ (.A1(_1128_),
    .A2(_0450_),
    .B1(_0571_),
    .B2(_0454_),
    .Y(_2072_));
 sky130_fd_sc_hd__a221oi_1 _5375_ (.A1(_3009_),
    .A2(_0930_),
    .B1(_3013_),
    .B2(_0931_),
    .C1(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__o22ai_1 _5376_ (.A1(_0811_),
    .A2(_0464_),
    .B1(_1559_),
    .B2(_0467_),
    .Y(_2074_));
 sky130_fd_sc_hd__a221oi_1 _5377_ (.A1(_2828_),
    .A2(_0936_),
    .B1(_2846_),
    .B2(_0937_),
    .C1(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(_0438_),
    .B(_2886_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand2_1 _5379_ (.A(_0442_),
    .B(_0695_),
    .Y(_2077_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(_2076_),
    .B(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__a221oi_1 _5381_ (.A1(_2839_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_2908_),
    .C1(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__nand2_1 _5382_ (.A(_0421_),
    .B(_0379_),
    .Y(_2080_));
 sky130_fd_sc_hd__nand2_1 _5383_ (.A(_0425_),
    .B(_0649_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_1 _5384_ (.A(_2080_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__a221oi_1 _5385_ (.A1(_0415_),
    .A2(_0426_),
    .B1(_0418_),
    .B2(_0707_),
    .C1(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__and4_1 _5386_ (.A(_2073_),
    .B(_2075_),
    .C(_2079_),
    .D(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__o22ai_1 _5387_ (.A1(_0606_),
    .A2(_0908_),
    .B1(_0342_),
    .B2(_0909_),
    .Y(_2085_));
 sky130_fd_sc_hd__a221oi_1 _5388_ (.A1(_3114_),
    .A2(_0906_),
    .B1(_3127_),
    .B2(_0907_),
    .C1(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__o22ai_2 _5389_ (.A1(_1580_),
    .A2(_0502_),
    .B1(_0671_),
    .B2(_0915_),
    .Y(_2087_));
 sky130_fd_sc_hd__a221oi_4 _5390_ (.A1(_2808_),
    .A2(_0918_),
    .B1(_2810_),
    .B2(_0917_),
    .C1(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__o22ai_1 _5391_ (.A1(_3122_),
    .A2(_0483_),
    .B1(_0618_),
    .B2(_0487_),
    .Y(_2089_));
 sky130_fd_sc_hd__a221oi_1 _5392_ (.A1(_3030_),
    .A2(_0478_),
    .B1(_0422_),
    .B2(_0480_),
    .C1(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__o22ai_1 _5393_ (.A1(_0902_),
    .A2(_0922_),
    .B1(_1406_),
    .B2(_0923_),
    .Y(_2091_));
 sky130_fd_sc_hd__a221oi_1 _5394_ (.A1(_3134_),
    .A2(_0925_),
    .B1(_2971_),
    .B2(_0926_),
    .C1(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__and4_1 _5395_ (.A(_2086_),
    .B(_2088_),
    .C(_2090_),
    .D(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__and4_1 _5396_ (.A(_2056_),
    .B(_2071_),
    .C(_2084_),
    .D(_2093_),
    .X(_2094_));
 sky130_fd_sc_hd__a22o_1 _5397_ (.A1(_2854_),
    .A2(_0647_),
    .B1(_2857_),
    .B2(_0430_),
    .X(_2095_));
 sky130_fd_sc_hd__a221oi_1 _5398_ (.A1(_2788_),
    .A2(_0825_),
    .B1(_0330_),
    .B2(_0824_),
    .C1(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _5399_ (.A(_2838_),
    .B(_0334_),
    .Y(_2097_));
 sky130_fd_sc_hd__nand2_1 _5400_ (.A(_2845_),
    .B(_2794_),
    .Y(_2098_));
 sky130_fd_sc_hd__nand2_1 _5401_ (.A(_2097_),
    .B(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__a221oi_1 _5402_ (.A1(_2786_),
    .A2(_2827_),
    .B1(_2792_),
    .B2(_2832_),
    .C1(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__nand2_1 _5403_ (.A(_2879_),
    .B(_2806_),
    .Y(_2101_));
 sky130_fd_sc_hd__o21ai_1 _5404_ (.A1(_1461_),
    .A2(_2870_),
    .B1(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__a31oi_1 _5405_ (.A1(_2812_),
    .A2(_2860_),
    .A3(_2874_),
    .B1(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__nand2_1 _5406_ (.A(_2890_),
    .B(_2800_),
    .Y(_2104_));
 sky130_fd_sc_hd__nand2_1 _5407_ (.A(_2894_),
    .B(_0648_),
    .Y(_2105_));
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_2104_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__a221oi_1 _5409_ (.A1(_2885_),
    .A2(_2796_),
    .B1(_2888_),
    .B2(_3078_),
    .C1(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__and4_1 _5410_ (.A(_2096_),
    .B(_2100_),
    .C(_2103_),
    .D(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__o22ai_1 _5411_ (.A1(_0724_),
    .A2(_2911_),
    .B1(_3018_),
    .B2(_2916_),
    .Y(_2109_));
 sky130_fd_sc_hd__a221oi_1 _5412_ (.A1(_0384_),
    .A2(_2903_),
    .B1(_3050_),
    .B2(_2907_),
    .C1(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(_2925_),
    .B(_0591_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_1 _5414_ (.A(_2928_),
    .B(_0524_),
    .Y(_2112_));
 sky130_fd_sc_hd__nand2_1 _5415_ (.A(_2111_),
    .B(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__a221oi_1 _5416_ (.A1(_2920_),
    .A2(_2790_),
    .B1(_2923_),
    .B2(_0436_),
    .C1(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__nand2_1 _5417_ (.A(_2944_),
    .B(_2814_),
    .Y(_2115_));
 sky130_fd_sc_hd__nand2_1 _5418_ (.A(_2948_),
    .B(_0566_),
    .Y(_2116_));
 sky130_fd_sc_hd__nand2_1 _5419_ (.A(_2115_),
    .B(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__a221oi_1 _5420_ (.A1(_3002_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_0589_),
    .C1(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__nand2_1 _5421_ (.A(_2961_),
    .B(_2777_),
    .Y(_2119_));
 sky130_fd_sc_hd__nand2_1 _5422_ (.A(_2965_),
    .B(_2798_),
    .Y(_2120_));
 sky130_fd_sc_hd__nand2_1 _5423_ (.A(_2119_),
    .B(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__a221oi_1 _5424_ (.A1(_0326_),
    .A2(_2955_),
    .B1(_0745_),
    .B2(_2959_),
    .C1(_2121_),
    .Y(_2122_));
 sky130_fd_sc_hd__and4_1 _5425_ (.A(_2110_),
    .B(_2114_),
    .C(_2118_),
    .D(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__nand2_1 _5426_ (.A(_2986_),
    .B(_0623_),
    .Y(_2124_));
 sky130_fd_sc_hd__o21ai_1 _5427_ (.A1(_0543_),
    .A2(_2984_),
    .B1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__a221oi_1 _5428_ (.A1(_2987_),
    .A2(_2976_),
    .B1(_2956_),
    .B2(_2981_),
    .C1(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__or2_1 _5429_ (.A(_0880_),
    .B(_0858_),
    .X(_2127_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(_2997_),
    .B(_2912_),
    .Y(_2128_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_3001_),
    .B(_2891_),
    .Y(_2129_));
 sky130_fd_sc_hd__o2111a_1 _5432_ (.A1(_0452_),
    .A2(_2993_),
    .B1(_2127_),
    .C1(_2128_),
    .D1(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__o22ai_1 _5433_ (.A1(_0490_),
    .A2(_3016_),
    .B1(_0346_),
    .B2(_3022_),
    .Y(_2131_));
 sky130_fd_sc_hd__a221oi_2 _5434_ (.A1(_0768_),
    .A2(_3008_),
    .B1(_3092_),
    .B2(_3012_),
    .C1(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__nand2_1 _5435_ (.A(_3035_),
    .B(_0537_),
    .Y(_2133_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(_3039_),
    .B(_0410_),
    .Y(_2134_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_2133_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__a221oi_1 _5438_ (.A1(_3028_),
    .A2(_3104_),
    .B1(_0631_),
    .B2(_3033_),
    .C1(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__and4_1 _5439_ (.A(_2126_),
    .B(_2130_),
    .C(_2132_),
    .D(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(_3052_),
    .B(_0391_),
    .Y(_2138_));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(_3057_),
    .B(_0395_),
    .Y(_2139_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_2138_),
    .B(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__a221oi_1 _5443_ (.A1(_3079_),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_3058_),
    .C1(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__nand2_1 _5444_ (.A(_3069_),
    .B(_2998_),
    .Y(_2142_));
 sky130_fd_sc_hd__nand2_1 _5445_ (.A(_3072_),
    .B(_0596_),
    .Y(_2143_));
 sky130_fd_sc_hd__nand2_1 _5446_ (.A(_2142_),
    .B(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__a221oi_1 _5447_ (.A1(_3063_),
    .A2(_0439_),
    .B1(_3066_),
    .B2(_2932_),
    .C1(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(_3088_),
    .B(_0459_),
    .Y(_2146_));
 sky130_fd_sc_hd__o21ai_1 _5449_ (.A1(_0795_),
    .A2(_3086_),
    .B1(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__a221oi_1 _5450_ (.A1(_3077_),
    .A2(_0457_),
    .B1(_0622_),
    .B2(_3082_),
    .C1(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__nand2_1 _5451_ (.A(_3100_),
    .B(_0471_),
    .Y(_2149_));
 sky130_fd_sc_hd__nand2_1 _5452_ (.A(_3103_),
    .B(_2865_),
    .Y(_2150_));
 sky130_fd_sc_hd__nand2_1 _5453_ (.A(_2149_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__a221oi_2 _5454_ (.A1(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0651_),
    .C1(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__and4_1 _5455_ (.A(_2141_),
    .B(_2145_),
    .C(_2148_),
    .D(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__and4_1 _5456_ (.A(_2108_),
    .B(_2123_),
    .C(_2137_),
    .D(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__nand3_2 _5457_ (.A(_2094_),
    .B(_2154_),
    .C(_3113_),
    .Y(_2155_));
 sky130_fd_sc_hd__o21a_1 _5458_ (.A1(_3083_),
    .A2(_0525_),
    .B1(_2776_),
    .X(_2156_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_2155_),
    .B(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__o21ai_1 _5460_ (.A1(_2776_),
    .A2(_2042_),
    .B1(_2157_),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _5461_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2158_));
 sky130_fd_sc_hd__a22o_1 _5462_ (.A1(_0426_),
    .A2(_0401_),
    .B1(_0404_),
    .B2(_0707_),
    .X(_2159_));
 sky130_fd_sc_hd__a221oi_1 _5463_ (.A1(_2817_),
    .A2(_0407_),
    .B1(_2865_),
    .B2(_0409_),
    .C1(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__nand2_1 _5464_ (.A(_0372_),
    .B(_0443_),
    .Y(_2161_));
 sky130_fd_sc_hd__o21ai_1 _5465_ (.A1(_0660_),
    .A2(_0369_),
    .B1(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__a221oi_2 _5466_ (.A1(_0651_),
    .A2(_0375_),
    .B1(_2828_),
    .B2(_0378_),
    .C1(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(_0390_),
    .B(_0622_),
    .Y(_2164_));
 sky130_fd_sc_hd__nand2_1 _5468_ (.A(_0394_),
    .B(_0422_),
    .Y(_2165_));
 sky130_fd_sc_hd__nand2_1 _5469_ (.A(_2164_),
    .B(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__a221oi_1 _5470_ (.A1(_0383_),
    .A2(_3058_),
    .B1(_3064_),
    .B2(_0388_),
    .C1(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__nand2_1 _5471_ (.A(_0360_),
    .B(_0323_),
    .Y(_2168_));
 sky130_fd_sc_hd__nand2_1 _5472_ (.A(_0363_),
    .B(_0352_),
    .Y(_2169_));
 sky130_fd_sc_hd__nand2_1 _5473_ (.A(_2168_),
    .B(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__a221oi_1 _5474_ (.A1(_0410_),
    .A2(_0355_),
    .B1(_0357_),
    .B2(_3114_),
    .C1(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__and4_1 _5475_ (.A(_2160_),
    .B(_2163_),
    .C(_2167_),
    .D(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__nor2_1 _5476_ (.A(_0902_),
    .B(_0347_),
    .Y(_2173_));
 sky130_fd_sc_hd__a31o_1 _5477_ (.A1(_0419_),
    .A2(_3055_),
    .A3(_2842_),
    .B1(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__a221oi_1 _5478_ (.A1(_3053_),
    .A2(_0341_),
    .B1(_3044_),
    .B2(_0337_),
    .C1(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__or2_1 _5479_ (.A(_0655_),
    .B(_3137_),
    .X(_2176_));
 sky130_fd_sc_hd__or2_1 _5480_ (.A(_0933_),
    .B(_3141_),
    .X(_2177_));
 sky130_fd_sc_hd__nand2_1 _5481_ (.A(_3144_),
    .B(_3067_),
    .Y(_2178_));
 sky130_fd_sc_hd__o2111a_1 _5482_ (.A1(_1880_),
    .A2(_3133_),
    .B1(_2176_),
    .C1(_2177_),
    .D1(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_0325_),
    .B(_0345_),
    .Y(_2180_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_0329_),
    .B(_0447_),
    .Y(_2181_));
 sky130_fd_sc_hd__nand2_1 _5485_ (.A(_2180_),
    .B(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__a221oi_2 _5486_ (.A1(_0484_),
    .A2(_3150_),
    .B1(_0322_),
    .B2(_0596_),
    .C1(_2182_),
    .Y(_2183_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(_3125_),
    .B(_0634_),
    .Y(_2184_));
 sky130_fd_sc_hd__o21ai_1 _5488_ (.A1(_2068_),
    .A2(_3123_),
    .B1(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__a221oi_2 _5489_ (.A1(_0385_),
    .A2(_3116_),
    .B1(_0613_),
    .B2(_3120_),
    .C1(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__and4_1 _5490_ (.A(_2175_),
    .B(_2179_),
    .C(_2183_),
    .D(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__o22ai_1 _5491_ (.A1(_1249_),
    .A2(_0450_),
    .B1(_0725_),
    .B2(_0454_),
    .Y(_2188_));
 sky130_fd_sc_hd__a221oi_1 _5492_ (.A1(_3013_),
    .A2(_0930_),
    .B1(_2956_),
    .B2(_0931_),
    .C1(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__o22ai_1 _5493_ (.A1(_0914_),
    .A2(_0464_),
    .B1(_1677_),
    .B2(_0467_),
    .Y(_2190_));
 sky130_fd_sc_hd__a221oi_1 _5494_ (.A1(_2846_),
    .A2(_0936_),
    .B1(_2886_),
    .B2(_0937_),
    .C1(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__nand2_1 _5495_ (.A(_0438_),
    .B(_2966_),
    .Y(_2192_));
 sky130_fd_sc_hd__nand2_1 _5496_ (.A(_0442_),
    .B(_2880_),
    .Y(_2193_));
 sky130_fd_sc_hd__nand2_1 _5497_ (.A(_2192_),
    .B(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__a221oi_1 _5498_ (.A1(_2899_),
    .A2(_0433_),
    .B1(_0435_),
    .B2(_2952_),
    .C1(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_0421_),
    .B(_0631_),
    .Y(_2196_));
 sky130_fd_sc_hd__nand2_1 _5500_ (.A(_0425_),
    .B(_3002_),
    .Y(_2197_));
 sky130_fd_sc_hd__nand2_1 _5501_ (.A(_2196_),
    .B(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__a221oi_1 _5502_ (.A1(_0415_),
    .A2(_2932_),
    .B1(_0418_),
    .B2(_3098_),
    .C1(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hd__and4_1 _5503_ (.A(_2189_),
    .B(_2191_),
    .C(_2195_),
    .D(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__o22ai_1 _5504_ (.A1(_3122_),
    .A2(_0908_),
    .B1(_0618_),
    .B2(_0909_),
    .Y(_2201_));
 sky130_fd_sc_hd__a221oi_1 _5505_ (.A1(_3127_),
    .A2(_0906_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .B2(_0907_),
    .C1(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__o22ai_2 _5506_ (.A1(_1698_),
    .A2(_0502_),
    .B1(_0811_),
    .B2(_0915_),
    .Y(_2203_));
 sky130_fd_sc_hd__a221oi_4 _5507_ (.A1(_2810_),
    .A2(_0918_),
    .B1(_2812_),
    .B2(_0917_),
    .C1(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__o22ai_1 _5508_ (.A1(_0342_),
    .A2(_0483_),
    .B1(_0764_),
    .B2(_0487_),
    .Y(_2205_));
 sky130_fd_sc_hd__a221oi_1 _5509_ (.A1(_0574_),
    .A2(_0478_),
    .B1(_3030_),
    .B2(_0480_),
    .C1(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__o22ai_1 _5510_ (.A1(_1043_),
    .A2(_0922_),
    .B1(_1527_),
    .B2(_0923_),
    .Y(_2207_));
 sky130_fd_sc_hd__a221oi_1 _5511_ (.A1(_2971_),
    .A2(_0925_),
    .B1(_3083_),
    .B2(_0926_),
    .C1(_2207_),
    .Y(_2208_));
 sky130_fd_sc_hd__and4_1 _5512_ (.A(_2202_),
    .B(_2204_),
    .C(_2206_),
    .D(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__and4_1 _5513_ (.A(_2172_),
    .B(_2187_),
    .C(_2200_),
    .D(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__a22o_1 _5514_ (.A1(_2854_),
    .A2(_0330_),
    .B1(_2857_),
    .B2(_0647_),
    .X(_2211_));
 sky130_fd_sc_hd__a221oi_1 _5515_ (.A1(_2790_),
    .A2(_0825_),
    .B1(_3134_),
    .B2(_0824_),
    .C1(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__nand2_1 _5516_ (.A(_2838_),
    .B(_0384_),
    .Y(_2213_));
 sky130_fd_sc_hd__nand2_1 _5517_ (.A(_2845_),
    .B(_2796_),
    .Y(_2214_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(_2213_),
    .B(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__a221oi_1 _5519_ (.A1(_2788_),
    .A2(_2827_),
    .B1(_2794_),
    .B2(_2832_),
    .C1(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__nand2_1 _5520_ (.A(_2878_),
    .B(_2808_),
    .Y(_2217_));
 sky130_fd_sc_hd__o21ai_1 _5521_ (.A1(_1580_),
    .A2(_2870_),
    .B1(_2217_),
    .Y(_2218_));
 sky130_fd_sc_hd__a31oi_1 _5522_ (.A1(_2814_),
    .A2(_2860_),
    .A3(_2874_),
    .B1(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(_2890_),
    .B(_2802_),
    .Y(_2220_));
 sky130_fd_sc_hd__nand2_1 _5524_ (.A(_2894_),
    .B(_2998_),
    .Y(_2221_));
 sky130_fd_sc_hd__nand2_1 _5525_ (.A(_2220_),
    .B(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__a221oi_1 _5526_ (.A1(_2885_),
    .A2(_2798_),
    .B1(_2888_),
    .B2(_0589_),
    .C1(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__and4_1 _5527_ (.A(_2212_),
    .B(_2216_),
    .C(_2219_),
    .D(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__o22ai_1 _5528_ (.A1(_0863_),
    .A2(_2911_),
    .B1(_0571_),
    .B2(_2916_),
    .Y(_2225_));
 sky130_fd_sc_hd__a221oi_1 _5529_ (.A1(_3050_),
    .A2(_2903_),
    .B1(_0358_),
    .B2(_2907_),
    .C1(_2225_),
    .Y(_2226_));
 sky130_fd_sc_hd__nand2_1 _5530_ (.A(_2925_),
    .B(_0436_),
    .Y(_2227_));
 sky130_fd_sc_hd__nand2_1 _5531_ (.A(_2928_),
    .B(_3078_),
    .Y(_2228_));
 sky130_fd_sc_hd__nand2_1 _5532_ (.A(_2227_),
    .B(_2228_),
    .Y(_2229_));
 sky130_fd_sc_hd__a221oi_1 _5533_ (.A1(_2920_),
    .A2(_2792_),
    .B1(_2923_),
    .B2(_0648_),
    .C1(_2229_),
    .Y(_2230_));
 sky130_fd_sc_hd__nand2_1 _5534_ (.A(_2944_),
    .B(_0524_),
    .Y(_2231_));
 sky130_fd_sc_hd__nand2_1 _5535_ (.A(_2948_),
    .B(_0430_),
    .Y(_2232_));
 sky130_fd_sc_hd__nand2_1 _5536_ (.A(_2231_),
    .B(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__a221oi_1 _5537_ (.A1(_3036_),
    .A2(_2939_),
    .B1(_2941_),
    .B2(_0591_),
    .C1(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__nand2_1 _5538_ (.A(_2961_),
    .B(_2786_),
    .Y(_2235_));
 sky130_fd_sc_hd__nand2_1 _5539_ (.A(_2965_),
    .B(_2800_),
    .Y(_2236_));
 sky130_fd_sc_hd__nand2_1 _5540_ (.A(_2235_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__a221oi_1 _5541_ (.A1(_3017_),
    .A2(_2955_),
    .B1(_0884_),
    .B2(_2959_),
    .C1(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__and4_1 _5542_ (.A(_2226_),
    .B(_2230_),
    .C(_2234_),
    .D(_2238_),
    .X(_2239_));
 sky130_fd_sc_hd__nand2_1 _5543_ (.A(_2986_),
    .B(_0768_),
    .Y(_2240_));
 sky130_fd_sc_hd__o21ai_1 _5544_ (.A1(_2913_),
    .A2(_2984_),
    .B1(_2240_),
    .Y(_2241_));
 sky130_fd_sc_hd__a221oi_1 _5545_ (.A1(_3005_),
    .A2(_2976_),
    .B1(_3147_),
    .B2(_2981_),
    .C1(_2241_),
    .Y(_2242_));
 sky130_fd_sc_hd__or2_1 _5546_ (.A(_2909_),
    .B(_0858_),
    .X(_2243_));
 sky130_fd_sc_hd__nand2_1 _5547_ (.A(_2997_),
    .B(_0451_),
    .Y(_2244_));
 sky130_fd_sc_hd__nand2_1 _5548_ (.A(_3001_),
    .B(_0537_),
    .Y(_2245_));
 sky130_fd_sc_hd__o2111a_1 _5549_ (.A1(_0656_),
    .A2(_2993_),
    .B1(_2243_),
    .C1(_2244_),
    .D1(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__o22ai_1 _5550_ (.A1(_0481_),
    .A2(_3016_),
    .B1(_0511_),
    .B2(_3022_),
    .Y(_2247_));
 sky130_fd_sc_hd__a221oi_2 _5551_ (.A1(_3092_),
    .A2(_3008_),
    .B1(_0595_),
    .B2(_3012_),
    .C1(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__nand2_1 _5552_ (.A(_3035_),
    .B(_0695_),
    .Y(_2249_));
 sky130_fd_sc_hd__nand2_1 _5553_ (.A(_3039_),
    .B(_3104_),
    .Y(_2250_));
 sky130_fd_sc_hd__nand2_1 _5554_ (.A(_2249_),
    .B(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__a221oi_1 _5555_ (.A1(_3028_),
    .A2(_0379_),
    .B1(_0471_),
    .B2(_3033_),
    .C1(_2251_),
    .Y(_2252_));
 sky130_fd_sc_hd__and4_1 _5556_ (.A(_2242_),
    .B(_2246_),
    .C(_2248_),
    .D(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__nand2_1 _5557_ (.A(_3052_),
    .B(_3079_),
    .Y(_2254_));
 sky130_fd_sc_hd__nand2_1 _5558_ (.A(_3057_),
    .B(_0479_),
    .Y(_2255_));
 sky130_fd_sc_hd__nand2_1 _5559_ (.A(_2254_),
    .B(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__a221oi_2 _5560_ (.A1(_0395_),
    .A2(_3047_),
    .B1(_3049_),
    .B2(_0513_),
    .C1(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__nand2_1 _5561_ (.A(_3069_),
    .B(_0566_),
    .Y(_2258_));
 sky130_fd_sc_hd__nand2_1 _5562_ (.A(_3072_),
    .B(_0746_),
    .Y(_2259_));
 sky130_fd_sc_hd__nand2_1 _5563_ (.A(_2258_),
    .B(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__a221oi_1 _5564_ (.A1(_3063_),
    .A2(_0649_),
    .B1(_3066_),
    .B2(_0550_),
    .C1(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__nand2_1 _5565_ (.A(_3088_),
    .B(_2977_),
    .Y(_2262_));
 sky130_fd_sc_hd__o21ai_1 _5566_ (.A1(_0932_),
    .A2(_3086_),
    .B1(_2262_),
    .Y(_2263_));
 sky130_fd_sc_hd__a221oi_1 _5567_ (.A1(_3077_),
    .A2(_0459_),
    .B1(_3029_),
    .B2(_3082_),
    .C1(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__nand2_1 _5568_ (.A(_3100_),
    .B(_0439_),
    .Y(_2265_));
 sky130_fd_sc_hd__nand2_1 _5569_ (.A(_3103_),
    .B(_2921_),
    .Y(_2266_));
 sky130_fd_sc_hd__nand2_1 _5570_ (.A(_2265_),
    .B(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__a221oi_1 _5571_ (.A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .A2(_3095_),
    .B1(_3097_),
    .B2(_0791_),
    .C1(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__and4_1 _5572_ (.A(_2257_),
    .B(_2261_),
    .C(_2264_),
    .D(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__and4_1 _5573_ (.A(_2224_),
    .B(_2239_),
    .C(_2253_),
    .D(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__nand3_1 _5574_ (.A(_2210_),
    .B(_2270_),
    .C(_3113_),
    .Y(_2271_));
 sky130_fd_sc_hd__o21a_1 _5575_ (.A1(_0457_),
    .A2(_0525_),
    .B1(_2776_),
    .X(_2272_));
 sky130_fd_sc_hd__nand2_1 _5576_ (.A(_2271_),
    .B(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__o21ai_1 _5577_ (.A1(_2776_),
    .A2(_2158_),
    .B1(_2273_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_4 _5578_ (.A(_2779_),
    .B(_2762_),
    .Y(_2274_));
 sky130_fd_sc_hd__buf_4 _5579_ (.A(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(net7),
    .A1(_0524_),
    .S(_2275_),
    .X(_2276_));
 sky130_fd_sc_hd__clkbuf_1 _5581_ (.A(_2276_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(net6),
    .A1(_3078_),
    .S(_2275_),
    .X(_2277_));
 sky130_fd_sc_hd__clkbuf_1 _5583_ (.A(_2277_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5584_ (.A0(net5),
    .A1(_0589_),
    .S(_2275_),
    .X(_2278_));
 sky130_fd_sc_hd__clkbuf_1 _5585_ (.A(_2278_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(net4),
    .A1(_0591_),
    .S(_2275_),
    .X(_2279_));
 sky130_fd_sc_hd__clkbuf_1 _5587_ (.A(_2279_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5588_ (.A0(net3),
    .A1(_0436_),
    .S(_2275_),
    .X(_2280_));
 sky130_fd_sc_hd__clkbuf_1 _5589_ (.A(_2280_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5590_ (.A0(net2),
    .A1(_0648_),
    .S(_2275_),
    .X(_2281_));
 sky130_fd_sc_hd__clkbuf_1 _5591_ (.A(_2281_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5592_ (.A0(net16),
    .A1(_2998_),
    .S(_2275_),
    .X(_2282_));
 sky130_fd_sc_hd__clkbuf_1 _5593_ (.A(_2282_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(net15),
    .A1(_0566_),
    .S(_2275_),
    .X(_2283_));
 sky130_fd_sc_hd__clkbuf_1 _5595_ (.A(_2283_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5596_ (.A0(net14),
    .A1(_0430_),
    .S(_2275_),
    .X(_2284_));
 sky130_fd_sc_hd__clkbuf_1 _5597_ (.A(_2284_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(net13),
    .A1(_0647_),
    .S(_2275_),
    .X(_2285_));
 sky130_fd_sc_hd__clkbuf_1 _5599_ (.A(_2285_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(net12),
    .A1(_0330_),
    .S(_2275_),
    .X(_2286_));
 sky130_fd_sc_hd__clkbuf_1 _5601_ (.A(_2286_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5602_ (.A0(net11),
    .A1(_3134_),
    .S(_2275_),
    .X(_2287_));
 sky130_fd_sc_hd__clkbuf_1 _5603_ (.A(_2287_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5604_ (.A0(net10),
    .A1(_2971_),
    .S(_2274_),
    .X(_2288_));
 sky130_fd_sc_hd__clkbuf_1 _5605_ (.A(_2288_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5606_ (.A0(net9),
    .A1(_3083_),
    .S(_2274_),
    .X(_2289_));
 sky130_fd_sc_hd__clkbuf_1 _5607_ (.A(_2289_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5608_ (.A0(net8),
    .A1(_0457_),
    .S(_2274_),
    .X(_2290_));
 sky130_fd_sc_hd__clkbuf_1 _5609_ (.A(_2290_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(net1),
    .A1(_0459_),
    .S(_2274_),
    .X(_2291_));
 sky130_fd_sc_hd__clkbuf_1 _5611_ (.A(_2291_),
    .X(_0267_));
 sky130_fd_sc_hd__or4b_4 _5612_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(_2761_),
    .D_N(_2779_),
    .X(_2292_));
 sky130_fd_sc_hd__buf_4 _5613_ (.A(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(net7),
    .A1(_2977_),
    .S(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__clkbuf_1 _5615_ (.A(_2294_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(net6),
    .A1(_2908_),
    .S(_2293_),
    .X(_2295_));
 sky130_fd_sc_hd__clkbuf_1 _5617_ (.A(_2295_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5618_ (.A0(net5),
    .A1(_2952_),
    .S(_2293_),
    .X(_2296_));
 sky130_fd_sc_hd__clkbuf_1 _5619_ (.A(_2296_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5620_ (.A0(net4),
    .A1(_2912_),
    .S(_2293_),
    .X(_2297_));
 sky130_fd_sc_hd__clkbuf_1 _5621_ (.A(_2297_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5622_ (.A0(net3),
    .A1(_0451_),
    .S(_2293_),
    .X(_2298_));
 sky130_fd_sc_hd__clkbuf_1 _5623_ (.A(_2298_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5624_ (.A0(net2),
    .A1(_2839_),
    .S(_2293_),
    .X(_2299_));
 sky130_fd_sc_hd__clkbuf_1 _5625_ (.A(_2299_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5626_ (.A0(net16),
    .A1(_2899_),
    .S(_2293_),
    .X(_2300_));
 sky130_fd_sc_hd__clkbuf_1 _5627_ (.A(_2300_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5628_ (.A0(net15),
    .A1(_2904_),
    .S(_2293_),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _5629_ (.A(_2301_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5630_ (.A0(net14),
    .A1(_0447_),
    .S(_2293_),
    .X(_2302_));
 sky130_fd_sc_hd__clkbuf_1 _5631_ (.A(_2302_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5632_ (.A0(net13),
    .A1(_2987_),
    .S(_2293_),
    .X(_2303_));
 sky130_fd_sc_hd__clkbuf_1 _5633_ (.A(_2303_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5634_ (.A0(net12),
    .A1(_3005_),
    .S(_2293_),
    .X(_2304_));
 sky130_fd_sc_hd__clkbuf_1 _5635_ (.A(_2304_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(net11),
    .A1(_3009_),
    .S(_2293_),
    .X(_2305_));
 sky130_fd_sc_hd__clkbuf_1 _5637_ (.A(_2305_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5638_ (.A0(net10),
    .A1(_3013_),
    .S(_2292_),
    .X(_2306_));
 sky130_fd_sc_hd__clkbuf_1 _5639_ (.A(_2306_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5640_ (.A0(net9),
    .A1(_2956_),
    .S(_2292_),
    .X(_2307_));
 sky130_fd_sc_hd__clkbuf_1 _5641_ (.A(_2307_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5642_ (.A0(net8),
    .A1(_3147_),
    .S(_2292_),
    .X(_2308_));
 sky130_fd_sc_hd__clkbuf_1 _5643_ (.A(_2308_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5644_ (.A0(net1),
    .A1(_0326_),
    .S(_2292_),
    .X(_2309_));
 sky130_fd_sc_hd__clkbuf_1 _5645_ (.A(_2309_),
    .X(_0251_));
 sky130_fd_sc_hd__or4b_4 _5646_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(_2760_),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .D_N(_2779_),
    .X(_2310_));
 sky130_fd_sc_hd__clkbuf_8 _5647_ (.A(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__mux2_1 _5648_ (.A0(net7),
    .A1(_3017_),
    .S(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__clkbuf_1 _5649_ (.A(_2312_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5650_ (.A0(net6),
    .A1(_0338_),
    .S(_2311_),
    .X(_2313_));
 sky130_fd_sc_hd__clkbuf_1 _5651_ (.A(_2313_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5652_ (.A0(net5),
    .A1(_0334_),
    .S(_2311_),
    .X(_2314_));
 sky130_fd_sc_hd__clkbuf_1 _5653_ (.A(_2314_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(net4),
    .A1(_0384_),
    .S(_2311_),
    .X(_2315_));
 sky130_fd_sc_hd__clkbuf_1 _5655_ (.A(_2315_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5656_ (.A0(net3),
    .A1(_3050_),
    .S(_2311_),
    .X(_2316_));
 sky130_fd_sc_hd__clkbuf_1 _5657_ (.A(_2316_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5658_ (.A0(net2),
    .A1(_0358_),
    .S(_2311_),
    .X(_2317_));
 sky130_fd_sc_hd__clkbuf_1 _5659_ (.A(_2317_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5660_ (.A0(net16),
    .A1(_0623_),
    .S(_2311_),
    .X(_2318_));
 sky130_fd_sc_hd__clkbuf_1 _5661_ (.A(_2318_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5662_ (.A0(net15),
    .A1(_0768_),
    .S(_2311_),
    .X(_2319_));
 sky130_fd_sc_hd__clkbuf_1 _5663_ (.A(_2319_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5664_ (.A0(net14),
    .A1(_3092_),
    .S(_2311_),
    .X(_2320_));
 sky130_fd_sc_hd__clkbuf_1 _5665_ (.A(_2320_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5666_ (.A0(net13),
    .A1(_0595_),
    .S(_2311_),
    .X(_2321_));
 sky130_fd_sc_hd__clkbuf_1 _5667_ (.A(_2321_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5668_ (.A0(net12),
    .A1(_0745_),
    .S(_2311_),
    .X(_2322_));
 sky130_fd_sc_hd__clkbuf_1 _5669_ (.A(_2322_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5670_ (.A0(net11),
    .A1(_0884_),
    .S(_2311_),
    .X(_2323_));
 sky130_fd_sc_hd__clkbuf_1 _5671_ (.A(_2323_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(net10),
    .A1(_0484_),
    .S(_2310_),
    .X(_2324_));
 sky130_fd_sc_hd__clkbuf_1 _5673_ (.A(_2324_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(net9),
    .A1(_0345_),
    .S(_2310_),
    .X(_2325_));
 sky130_fd_sc_hd__clkbuf_1 _5675_ (.A(_2325_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(net8),
    .A1(_0510_),
    .S(_2310_),
    .X(_2326_));
 sky130_fd_sc_hd__clkbuf_1 _5677_ (.A(_2326_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(net1),
    .A1(_3053_),
    .S(_2310_),
    .X(_2327_));
 sky130_fd_sc_hd__clkbuf_1 _5679_ (.A(_2327_),
    .X(_0235_));
 sky130_fd_sc_hd__or2_4 _5680_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(_2781_),
    .X(_2328_));
 sky130_fd_sc_hd__buf_4 _5681_ (.A(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__mux2_1 _5682_ (.A0(net7),
    .A1(_3044_),
    .S(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__clkbuf_1 _5683_ (.A(_2330_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(net6),
    .A1(_3058_),
    .S(_2329_),
    .X(_2331_));
 sky130_fd_sc_hd__clkbuf_1 _5685_ (.A(_2331_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5686_ (.A0(net5),
    .A1(_0513_),
    .S(_2329_),
    .X(_2332_));
 sky130_fd_sc_hd__clkbuf_1 _5687_ (.A(_2332_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5688_ (.A0(net4),
    .A1(_3114_),
    .S(_2329_),
    .X(_2333_));
 sky130_fd_sc_hd__clkbuf_1 _5689_ (.A(_2333_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5690_ (.A0(net3),
    .A1(_3127_),
    .S(_2329_),
    .X(_2334_));
 sky130_fd_sc_hd__clkbuf_1 _5691_ (.A(_2334_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5692_ (.A0(net2),
    .A1(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .S(_2329_),
    .X(_2335_));
 sky130_fd_sc_hd__clkbuf_1 _5693_ (.A(_2335_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5694_ (.A0(net16),
    .A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .S(_2329_),
    .X(_2336_));
 sky130_fd_sc_hd__clkbuf_1 _5695_ (.A(_2336_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(net15),
    .A1(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .S(_2329_),
    .X(_2337_));
 sky130_fd_sc_hd__clkbuf_1 _5697_ (.A(_2337_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(net14),
    .A1(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .S(_2329_),
    .X(_2338_));
 sky130_fd_sc_hd__clkbuf_1 _5699_ (.A(_2338_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(net13),
    .A1(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .S(_2329_),
    .X(_2339_));
 sky130_fd_sc_hd__clkbuf_1 _5701_ (.A(_2339_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(net12),
    .A1(_3118_),
    .S(_2329_),
    .X(_2340_));
 sky130_fd_sc_hd__clkbuf_1 _5703_ (.A(_2340_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5704_ (.A0(net11),
    .A1(_0364_),
    .S(_2329_),
    .X(_2341_));
 sky130_fd_sc_hd__clkbuf_1 _5705_ (.A(_2341_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5706_ (.A0(net10),
    .A1(_0391_),
    .S(_2328_),
    .X(_2342_));
 sky130_fd_sc_hd__clkbuf_1 _5707_ (.A(_2342_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(net9),
    .A1(_3079_),
    .S(_2328_),
    .X(_2343_));
 sky130_fd_sc_hd__clkbuf_1 _5709_ (.A(_2343_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(net8),
    .A1(_0395_),
    .S(_2328_),
    .X(_2344_));
 sky130_fd_sc_hd__clkbuf_1 _5711_ (.A(_2344_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5712_ (.A0(net1),
    .A1(_0479_),
    .S(_2328_),
    .X(_2345_));
 sky130_fd_sc_hd__clkbuf_1 _5713_ (.A(_2345_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_2 _5714_ (.A(_2779_),
    .B(_2765_),
    .Y(_2346_));
 sky130_fd_sc_hd__buf_4 _5715_ (.A(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(net7),
    .A1(_0475_),
    .S(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__clkbuf_1 _5717_ (.A(_2348_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(net6),
    .A1(_0385_),
    .S(_2347_),
    .X(_2349_));
 sky130_fd_sc_hd__clkbuf_1 _5719_ (.A(_2349_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(net5),
    .A1(_0634_),
    .S(_2347_),
    .X(_2350_));
 sky130_fd_sc_hd__clkbuf_1 _5721_ (.A(_2350_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5722_ (.A0(net4),
    .A1(_0416_),
    .S(_2347_),
    .X(_2351_));
 sky130_fd_sc_hd__clkbuf_1 _5723_ (.A(_2351_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5724_ (.A0(net3),
    .A1(_3067_),
    .S(_2347_),
    .X(_2352_));
 sky130_fd_sc_hd__clkbuf_1 _5725_ (.A(_2352_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _5726_ (.A0(net2),
    .A1(_0584_),
    .S(_2347_),
    .X(_2353_));
 sky130_fd_sc_hd__clkbuf_1 _5727_ (.A(_2353_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5728_ (.A0(net16),
    .A1(_0419_),
    .S(_2347_),
    .X(_2354_));
 sky130_fd_sc_hd__clkbuf_1 _5729_ (.A(_2354_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _5730_ (.A0(net15),
    .A1(_0323_),
    .S(_2347_),
    .X(_2355_));
 sky130_fd_sc_hd__clkbuf_1 _5731_ (.A(_2355_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _5732_ (.A0(net14),
    .A1(_0613_),
    .S(_2347_),
    .X(_2356_));
 sky130_fd_sc_hd__clkbuf_1 _5733_ (.A(_2356_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(net13),
    .A1(_0352_),
    .S(_2347_),
    .X(_2357_));
 sky130_fd_sc_hd__clkbuf_1 _5735_ (.A(_2357_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _5736_ (.A0(net12),
    .A1(_0622_),
    .S(_2347_),
    .X(_2358_));
 sky130_fd_sc_hd__clkbuf_1 _5737_ (.A(_2358_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _5738_ (.A0(net11),
    .A1(_3029_),
    .S(_2347_),
    .X(_2359_));
 sky130_fd_sc_hd__clkbuf_1 _5739_ (.A(_2359_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _5740_ (.A0(net10),
    .A1(_0422_),
    .S(_2346_),
    .X(_2360_));
 sky130_fd_sc_hd__clkbuf_1 _5741_ (.A(_2360_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _5742_ (.A0(net9),
    .A1(_3030_),
    .S(_2346_),
    .X(_2361_));
 sky130_fd_sc_hd__clkbuf_1 _5743_ (.A(_2361_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(net8),
    .A1(_0574_),
    .S(_2346_),
    .X(_2362_));
 sky130_fd_sc_hd__clkbuf_1 _5745_ (.A(_2362_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _5746_ (.A0(net1),
    .A1(_3064_),
    .S(_2346_),
    .X(_2363_));
 sky130_fd_sc_hd__clkbuf_1 _5747_ (.A(_2363_),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(_2781_),
    .B(_2759_),
    .Y(_2364_));
 sky130_fd_sc_hd__and2_1 _5749_ (.A(_2784_),
    .B(_2364_),
    .X(_2365_));
 sky130_fd_sc_hd__clkbuf_1 _5750_ (.A(_2365_),
    .X(_0202_));
 sky130_fd_sc_hd__nand2_1 _5751_ (.A(_2780_),
    .B(_2760_),
    .Y(_2366_));
 sky130_fd_sc_hd__and2_1 _5752_ (.A(_2781_),
    .B(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__clkbuf_1 _5753_ (.A(_2367_),
    .X(_0201_));
 sky130_fd_sc_hd__or2_1 _5754_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .B(_2779_),
    .X(_2368_));
 sky130_fd_sc_hd__and2_1 _5755_ (.A(_2368_),
    .B(_2780_),
    .X(_2369_));
 sky130_fd_sc_hd__clkbuf_1 _5756_ (.A(_2369_),
    .X(_0200_));
 sky130_fd_sc_hd__or4b_4 _5757_ (.A(_2759_),
    .B(_2760_),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .D_N(_2779_),
    .X(_2370_));
 sky130_fd_sc_hd__buf_4 _5758_ (.A(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(net7),
    .A1(_0443_),
    .S(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__clkbuf_1 _5760_ (.A(_2372_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5761_ (.A0(net6),
    .A1(_0651_),
    .S(_2371_),
    .X(_2373_));
 sky130_fd_sc_hd__clkbuf_1 _5762_ (.A(_2373_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _5763_ (.A0(net5),
    .A1(_0791_),
    .S(_2371_),
    .X(_2374_));
 sky130_fd_sc_hd__clkbuf_1 _5764_ (.A(_2374_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(net4),
    .A1(_2962_),
    .S(_2371_),
    .X(_2375_));
 sky130_fd_sc_hd__clkbuf_1 _5766_ (.A(_2375_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _5767_ (.A0(net3),
    .A1(_2817_),
    .S(_2371_),
    .X(_2376_));
 sky130_fd_sc_hd__clkbuf_1 _5768_ (.A(_2376_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _5769_ (.A0(net2),
    .A1(_2865_),
    .S(_2371_),
    .X(_2377_));
 sky130_fd_sc_hd__clkbuf_1 _5770_ (.A(_2377_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(net16),
    .A1(_2921_),
    .S(_2371_),
    .X(_2378_));
 sky130_fd_sc_hd__clkbuf_1 _5772_ (.A(_2378_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _5773_ (.A0(net15),
    .A1(_2828_),
    .S(_2371_),
    .X(_2379_));
 sky130_fd_sc_hd__clkbuf_1 _5774_ (.A(_2379_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _5775_ (.A0(net14),
    .A1(_2846_),
    .S(_2371_),
    .X(_2380_));
 sky130_fd_sc_hd__clkbuf_1 _5776_ (.A(_2380_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _5777_ (.A0(net13),
    .A1(_2886_),
    .S(_2371_),
    .X(_2381_));
 sky130_fd_sc_hd__clkbuf_1 _5778_ (.A(_2381_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(net12),
    .A1(_2966_),
    .S(_2371_),
    .X(_2382_));
 sky130_fd_sc_hd__clkbuf_1 _5780_ (.A(_2382_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(net11),
    .A1(_2891_),
    .S(_2371_),
    .X(_2383_));
 sky130_fd_sc_hd__clkbuf_1 _5782_ (.A(_2383_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(net10),
    .A1(_0537_),
    .S(_2370_),
    .X(_2384_));
 sky130_fd_sc_hd__clkbuf_1 _5784_ (.A(_2384_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(net9),
    .A1(_0695_),
    .S(_2370_),
    .X(_2385_));
 sky130_fd_sc_hd__clkbuf_1 _5786_ (.A(_2385_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(net8),
    .A1(_2880_),
    .S(_2370_),
    .X(_2386_));
 sky130_fd_sc_hd__clkbuf_1 _5788_ (.A(_2386_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(net1),
    .A1(_0507_),
    .S(_2370_),
    .X(_2387_));
 sky130_fd_sc_hd__clkbuf_1 _5790_ (.A(_2387_),
    .X(_0184_));
 sky130_fd_sc_hd__or4b_4 _5791_ (.A(_2759_),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(_2761_),
    .D_N(_2779_),
    .X(_2388_));
 sky130_fd_sc_hd__buf_4 _5792_ (.A(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(net7),
    .A1(_0426_),
    .S(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_1 _5794_ (.A(_2390_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5795_ (.A0(net6),
    .A1(_2932_),
    .S(_2389_),
    .X(_2391_));
 sky130_fd_sc_hd__clkbuf_1 _5796_ (.A(_2391_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(net5),
    .A1(_0550_),
    .S(_2389_),
    .X(_2392_));
 sky130_fd_sc_hd__clkbuf_1 _5798_ (.A(_2392_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5799_ (.A0(net4),
    .A1(_0707_),
    .S(_2389_),
    .X(_2393_));
 sky130_fd_sc_hd__clkbuf_1 _5800_ (.A(_2393_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _5801_ (.A0(net3),
    .A1(_3098_),
    .S(_2389_),
    .X(_2394_));
 sky130_fd_sc_hd__clkbuf_1 _5802_ (.A(_2394_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5803_ (.A0(net2),
    .A1(_0596_),
    .S(_2389_),
    .X(_2395_));
 sky130_fd_sc_hd__clkbuf_1 _5804_ (.A(_2395_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5805_ (.A0(net16),
    .A1(_0746_),
    .S(_2389_),
    .X(_2396_));
 sky130_fd_sc_hd__clkbuf_1 _5806_ (.A(_2396_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(net15),
    .A1(_0410_),
    .S(_2389_),
    .X(_2397_));
 sky130_fd_sc_hd__clkbuf_1 _5808_ (.A(_2397_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5809_ (.A0(net14),
    .A1(_3104_),
    .S(_2389_),
    .X(_2398_));
 sky130_fd_sc_hd__clkbuf_1 _5810_ (.A(_2398_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5811_ (.A0(net13),
    .A1(_0379_),
    .S(_2389_),
    .X(_2399_));
 sky130_fd_sc_hd__clkbuf_1 _5812_ (.A(_2399_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5813_ (.A0(net12),
    .A1(_0631_),
    .S(_2389_),
    .X(_2400_));
 sky130_fd_sc_hd__clkbuf_1 _5814_ (.A(_2400_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5815_ (.A0(net11),
    .A1(_0471_),
    .S(_2389_),
    .X(_2401_));
 sky130_fd_sc_hd__clkbuf_1 _5816_ (.A(_2401_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5817_ (.A0(net10),
    .A1(_0439_),
    .S(_2388_),
    .X(_2402_));
 sky130_fd_sc_hd__clkbuf_1 _5818_ (.A(_2402_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _5819_ (.A0(net9),
    .A1(_0649_),
    .S(_2388_),
    .X(_2403_));
 sky130_fd_sc_hd__clkbuf_1 _5820_ (.A(_2403_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5821_ (.A0(net8),
    .A1(_3002_),
    .S(_2388_),
    .X(_2404_));
 sky130_fd_sc_hd__clkbuf_1 _5822_ (.A(_2404_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5823_ (.A0(net1),
    .A1(_3036_),
    .S(_2388_),
    .X(_2405_));
 sky130_fd_sc_hd__clkbuf_1 _5824_ (.A(_2405_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(net17),
    .B(net18),
    .Y(_2406_));
 sky130_fd_sc_hd__inv_2 _5826_ (.A(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__and3b_1 _5827_ (.A_N(net21),
    .B(_2407_),
    .C(net20),
    .X(_2408_));
 sky130_fd_sc_hd__inv_2 _5828_ (.A(\egd_top.exp_golomb_decoding.te_range[2] ),
    .Y(_2409_));
 sky130_fd_sc_hd__and2_2 _5829_ (.A(_2408_),
    .B(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__nor2_1 _5830_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2411_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(_2411_),
    .B(_2775_),
    .Y(_2412_));
 sky130_fd_sc_hd__inv_2 _5832_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2413_));
 sky130_fd_sc_hd__inv_4 _5833_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2414_));
 sky130_fd_sc_hd__nand2_1 _5834_ (.A(_2413_),
    .B(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__nor2_1 _5835_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(_2415_),
    .Y(_2416_));
 sky130_fd_sc_hd__inv_2 _5836_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_2417_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_2416_),
    .B(_2417_),
    .Y(_2418_));
 sky130_fd_sc_hd__inv_2 _5838_ (.A(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__inv_2 _5839_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2420_));
 sky130_fd_sc_hd__inv_2 _5840_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_2421_));
 sky130_fd_sc_hd__and3_1 _5841_ (.A(_2419_),
    .B(_2420_),
    .C(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__inv_2 _5842_ (.A(_2422_),
    .Y(_2423_));
 sky130_fd_sc_hd__nor2_1 _5843_ (.A(_2412_),
    .B(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__nor2_1 _5844_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2425_));
 sky130_fd_sc_hd__inv_2 _5845_ (.A(_2425_),
    .Y(_2426_));
 sky130_fd_sc_hd__nor2_1 _5846_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2426_),
    .Y(_2427_));
 sky130_fd_sc_hd__inv_2 _5847_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2428_));
 sky130_fd_sc_hd__nand2_1 _5848_ (.A(_2427_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__inv_2 _5849_ (.A(_2412_),
    .Y(_2430_));
 sky130_fd_sc_hd__nor2_1 _5850_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2431_));
 sky130_fd_sc_hd__nand2_2 _5851_ (.A(_2430_),
    .B(_2431_),
    .Y(_2432_));
 sky130_fd_sc_hd__a21o_1 _5852_ (.A1(_2422_),
    .A2(_2429_),
    .B1(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__nor2_2 _5853_ (.A(_2424_),
    .B(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__inv_6 _5854_ (.A(_2434_),
    .Y(_2435_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_2042_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2436_));
 sky130_fd_sc_hd__nand2_1 _5856_ (.A(_2436_),
    .B(_1926_),
    .Y(_2437_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(_2437_),
    .B(_2428_),
    .Y(_2438_));
 sky130_fd_sc_hd__inv_2 _5858_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2439_));
 sky130_fd_sc_hd__nand2_1 _5859_ (.A(_2438_),
    .B(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__inv_2 _5860_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2441_));
 sky130_fd_sc_hd__nand2_1 _5861_ (.A(_2440_),
    .B(_2441_),
    .Y(_2442_));
 sky130_fd_sc_hd__inv_2 _5862_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2443_));
 sky130_fd_sc_hd__nand2_1 _5863_ (.A(_2442_),
    .B(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(_2444_),
    .B(_2421_),
    .Y(_2445_));
 sky130_fd_sc_hd__nand2_1 _5865_ (.A(_2445_),
    .B(_2420_),
    .Y(_2446_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(_2446_),
    .B(_2419_),
    .Y(_2447_));
 sky130_fd_sc_hd__a21oi_1 _5867_ (.A1(_2413_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2448_));
 sky130_fd_sc_hd__nand2_1 _5868_ (.A(_2447_),
    .B(_2448_),
    .Y(_2449_));
 sky130_fd_sc_hd__nand2_2 _5869_ (.A(_2449_),
    .B(_2411_),
    .Y(_2450_));
 sky130_fd_sc_hd__o21ai_1 _5870_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_2428_),
    .Y(_2451_));
 sky130_fd_sc_hd__o211a_1 _5871_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .A2(_2451_),
    .B1(_2443_),
    .C1(_2441_),
    .X(_2452_));
 sky130_fd_sc_hd__a21o_1 _5872_ (.A1(_2418_),
    .A2(_2431_),
    .B1(_2412_),
    .X(_2453_));
 sky130_fd_sc_hd__o21bai_4 _5873_ (.A1(_2452_),
    .A2(_2423_),
    .B1_N(_2453_),
    .Y(_2454_));
 sky130_fd_sc_hd__nor2_2 _5874_ (.A(_2816_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_2455_));
 sky130_fd_sc_hd__nand3_1 _5875_ (.A(_2450_),
    .B(_2454_),
    .C(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hd__nor2_1 _5876_ (.A(_2435_),
    .B(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__inv_2 _5877_ (.A(_2457_),
    .Y(_2458_));
 sky130_fd_sc_hd__nor2_1 _5878_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .B(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__inv_2 _5879_ (.A(_2454_),
    .Y(_2460_));
 sky130_fd_sc_hd__nor2_1 _5880_ (.A(_2460_),
    .B(_2435_),
    .Y(_2461_));
 sky130_fd_sc_hd__nand2_2 _5881_ (.A(_2450_),
    .B(_2455_),
    .Y(_2462_));
 sky130_fd_sc_hd__nand2_1 _5882_ (.A(_2461_),
    .B(_2462_),
    .Y(_2463_));
 sky130_fd_sc_hd__nand2_1 _5883_ (.A(_2460_),
    .B(_2432_),
    .Y(_2464_));
 sky130_fd_sc_hd__inv_2 _5884_ (.A(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__nand3_1 _5885_ (.A(_2465_),
    .B(_2462_),
    .C(_2414_),
    .Y(_2466_));
 sky130_fd_sc_hd__o21ai_1 _5886_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .A2(_2463_),
    .B1(_2466_),
    .Y(_2467_));
 sky130_fd_sc_hd__nor2_1 _5887_ (.A(_2459_),
    .B(_2467_),
    .Y(_2468_));
 sky130_fd_sc_hd__nand3_4 _5888_ (.A(_2450_),
    .B(_2460_),
    .C(_2455_),
    .Y(_2469_));
 sky130_fd_sc_hd__inv_2 _5889_ (.A(_2469_),
    .Y(_2470_));
 sky130_fd_sc_hd__and3_1 _5890_ (.A(_2470_),
    .B(_2420_),
    .C(_2432_),
    .X(_2471_));
 sky130_fd_sc_hd__inv_2 _5891_ (.A(_2456_),
    .Y(_2472_));
 sky130_fd_sc_hd__and3_1 _5892_ (.A(_2472_),
    .B(_0684_),
    .C(_2432_),
    .X(_2473_));
 sky130_fd_sc_hd__nor2_1 _5893_ (.A(_2471_),
    .B(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__o21ai_1 _5894_ (.A1(_2435_),
    .A2(_2469_),
    .B1(_1926_),
    .Y(_2475_));
 sky130_fd_sc_hd__nor2_4 _5895_ (.A(_2435_),
    .B(_2469_),
    .Y(_2476_));
 sky130_fd_sc_hd__nand2_1 _5896_ (.A(_2476_),
    .B(_2158_),
    .Y(_2477_));
 sky130_fd_sc_hd__nand2_2 _5897_ (.A(_2475_),
    .B(_2477_),
    .Y(_2478_));
 sky130_fd_sc_hd__nor2_2 _5898_ (.A(_2454_),
    .B(_2435_),
    .Y(_2479_));
 sky130_fd_sc_hd__nand2_1 _5899_ (.A(_2478_),
    .B(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__nand3_2 _5900_ (.A(_2468_),
    .B(_2474_),
    .C(_2480_),
    .Y(_2481_));
 sky130_fd_sc_hd__nand2_2 _5901_ (.A(_2481_),
    .B(_2749_),
    .Y(_2482_));
 sky130_fd_sc_hd__inv_2 _5902_ (.A(_2482_),
    .Y(_2483_));
 sky130_fd_sc_hd__or2_1 _5903_ (.A(_2410_),
    .B(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__inv_2 _5904_ (.A(_2749_),
    .Y(_2485_));
 sky130_fd_sc_hd__a311o_1 _5905_ (.A1(_2462_),
    .A2(_2433_),
    .A3(_2454_),
    .B1(_2485_),
    .C1(_2424_),
    .X(_2486_));
 sky130_fd_sc_hd__nand2_1 _5906_ (.A(_2486_),
    .B(_2410_),
    .Y(_2487_));
 sky130_fd_sc_hd__nor2_1 _5907_ (.A(net18),
    .B(_2745_),
    .Y(_2488_));
 sky130_fd_sc_hd__nand2_1 _5908_ (.A(_2470_),
    .B(_2434_),
    .Y(_2489_));
 sky130_fd_sc_hd__nand2_1 _5909_ (.A(_2489_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2490_));
 sky130_fd_sc_hd__nand2_1 _5910_ (.A(_2476_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2491_));
 sky130_fd_sc_hd__nand2_1 _5911_ (.A(_2490_),
    .B(_2491_),
    .Y(_2492_));
 sky130_fd_sc_hd__o21ai_1 _5912_ (.A1(_2435_),
    .A2(_2469_),
    .B1(_2428_),
    .Y(_2493_));
 sky130_fd_sc_hd__nand3_1 _5913_ (.A(_2470_),
    .B(_2042_),
    .C(_2434_),
    .Y(_2494_));
 sky130_fd_sc_hd__nand2_1 _5914_ (.A(_2493_),
    .B(_2494_),
    .Y(_2495_));
 sky130_fd_sc_hd__nand2_1 _5915_ (.A(_2492_),
    .B(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__o21ai_1 _5916_ (.A1(_2435_),
    .A2(_2469_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2497_));
 sky130_fd_sc_hd__nand3_1 _5917_ (.A(_2470_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .C(_2434_),
    .Y(_2498_));
 sky130_fd_sc_hd__nand2_1 _5918_ (.A(_2497_),
    .B(_2498_),
    .Y(_2499_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_2478_),
    .B(_2499_),
    .Y(_2500_));
 sky130_fd_sc_hd__nand3_1 _5920_ (.A(_2496_),
    .B(_2500_),
    .C(_2479_),
    .Y(_2501_));
 sky130_fd_sc_hd__and2_1 _5921_ (.A(_2470_),
    .B(_2432_),
    .X(_2502_));
 sky130_fd_sc_hd__nor2_1 _5922_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2503_));
 sky130_fd_sc_hd__inv_2 _5923_ (.A(_2503_),
    .Y(_2504_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2505_));
 sky130_fd_sc_hd__nand2_1 _5925_ (.A(_2504_),
    .B(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__nand2_1 _5926_ (.A(_2502_),
    .B(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__xnor2_1 _5927_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2508_));
 sky130_fd_sc_hd__nand3_1 _5928_ (.A(_2472_),
    .B(_2432_),
    .C(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__nand2_1 _5929_ (.A(_2507_),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__xor2_1 _5930_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .X(_2511_));
 sky130_fd_sc_hd__nand2_1 _5931_ (.A(_2465_),
    .B(_2462_),
    .Y(_2512_));
 sky130_fd_sc_hd__nor2_1 _5932_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2513_));
 sky130_fd_sc_hd__inv_2 _5933_ (.A(_2513_),
    .Y(_2514_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2515_));
 sky130_fd_sc_hd__nand2_1 _5935_ (.A(_2514_),
    .B(_2515_),
    .Y(_2516_));
 sky130_fd_sc_hd__nand3_1 _5936_ (.A(_2461_),
    .B(_2462_),
    .C(_2516_),
    .Y(_2517_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2518_));
 sky130_fd_sc_hd__nand2_1 _5938_ (.A(_2426_),
    .B(_2518_),
    .Y(_2519_));
 sky130_fd_sc_hd__nand2_1 _5939_ (.A(_2457_),
    .B(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__o211ai_1 _5940_ (.A1(_2511_),
    .A2(_2512_),
    .B1(_2517_),
    .C1(_2520_),
    .Y(_2521_));
 sky130_fd_sc_hd__nor2_1 _5941_ (.A(_2510_),
    .B(_2521_),
    .Y(_2522_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_2501_),
    .B(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__nand3_1 _5943_ (.A(_2523_),
    .B(_2749_),
    .C(_2481_),
    .Y(_2524_));
 sky130_fd_sc_hd__nor2_2 _5944_ (.A(net17),
    .B(_2746_),
    .Y(_2525_));
 sky130_fd_sc_hd__a22o_1 _5945_ (.A1(_2483_),
    .A2(_2488_),
    .B1(_2524_),
    .B2(_2525_),
    .X(_2526_));
 sky130_fd_sc_hd__nand2_2 _5946_ (.A(_2523_),
    .B(_2749_),
    .Y(_2527_));
 sky130_fd_sc_hd__nand2_1 _5947_ (.A(_2527_),
    .B(_2482_),
    .Y(_2528_));
 sky130_fd_sc_hd__a32o_1 _5948_ (.A1(_2407_),
    .A2(_2484_),
    .A3(_2487_),
    .B1(_2526_),
    .B2(_2528_),
    .X(net20));
 sky130_fd_sc_hd__a31o_1 _5949_ (.A1(_2408_),
    .A2(net18),
    .A3(_2409_),
    .B1(_2745_),
    .X(_2529_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_2478_),
    .B(_2495_),
    .Y(_2530_));
 sky130_fd_sc_hd__o21ai_1 _5951_ (.A1(_2435_),
    .A2(_2469_),
    .B1(_2439_),
    .Y(_2531_));
 sky130_fd_sc_hd__nand2_1 _5952_ (.A(_2476_),
    .B(_1926_),
    .Y(_2532_));
 sky130_fd_sc_hd__nand2_1 _5953_ (.A(_2531_),
    .B(_2532_),
    .Y(_2533_));
 sky130_fd_sc_hd__nand2_1 _5954_ (.A(_2530_),
    .B(_2533_),
    .Y(_2534_));
 sky130_fd_sc_hd__o21ai_1 _5955_ (.A1(_2435_),
    .A2(_2469_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2535_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_2476_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2536_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(_2535_),
    .B(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__nand3_1 _5958_ (.A(_2478_),
    .B(_2537_),
    .C(_2495_),
    .Y(_2538_));
 sky130_fd_sc_hd__nand3_1 _5959_ (.A(_2534_),
    .B(_2538_),
    .C(_2479_),
    .Y(_2539_));
 sky130_fd_sc_hd__nor2_1 _5960_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2504_),
    .Y(_2540_));
 sky130_fd_sc_hd__nor2_1 _5961_ (.A(_2414_),
    .B(_2503_),
    .Y(_2541_));
 sky130_fd_sc_hd__o21ai_1 _5962_ (.A1(_2540_),
    .A2(_2541_),
    .B1(_2502_),
    .Y(_2542_));
 sky130_fd_sc_hd__nor2_1 _5963_ (.A(_2443_),
    .B(_2425_),
    .Y(_2543_));
 sky130_fd_sc_hd__o21ai_1 _5964_ (.A1(_2427_),
    .A2(_2543_),
    .B1(_2457_),
    .Y(_2544_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_2542_),
    .B(_2544_),
    .Y(_2545_));
 sky130_fd_sc_hd__and2_1 _5966_ (.A(_2415_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .X(_2546_));
 sky130_fd_sc_hd__nor2_1 _5967_ (.A(_2416_),
    .B(_2546_),
    .Y(_2547_));
 sky130_fd_sc_hd__nor2_1 _5968_ (.A(_2420_),
    .B(_2513_),
    .Y(_2548_));
 sky130_fd_sc_hd__nor2_1 _5969_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2514_),
    .Y(_2549_));
 sky130_fd_sc_hd__inv_2 _5970_ (.A(_2463_),
    .Y(_2550_));
 sky130_fd_sc_hd__o21ai_1 _5971_ (.A1(_2548_),
    .A2(_2549_),
    .B1(_2550_),
    .Y(_2551_));
 sky130_fd_sc_hd__o21ai_1 _5972_ (.A1(_2512_),
    .A2(_2547_),
    .B1(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__nor2_1 _5973_ (.A(_2545_),
    .B(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__nand2_1 _5974_ (.A(_2539_),
    .B(_2553_),
    .Y(_2554_));
 sky130_fd_sc_hd__nand2_2 _5975_ (.A(_2554_),
    .B(_2749_),
    .Y(_2555_));
 sky130_fd_sc_hd__or2_1 _5976_ (.A(_2527_),
    .B(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__nand2_2 _5977_ (.A(_2555_),
    .B(_2527_),
    .Y(_2557_));
 sky130_fd_sc_hd__nand3_1 _5978_ (.A(_2556_),
    .B(_2557_),
    .C(_2525_),
    .Y(_2558_));
 sky130_fd_sc_hd__o21ai_2 _5979_ (.A1(_2527_),
    .A2(_2529_),
    .B1(_2558_),
    .Y(net21));
 sky130_fd_sc_hd__o21ai_1 _5980_ (.A1(_2527_),
    .A2(_2555_),
    .B1(_2483_),
    .Y(_2559_));
 sky130_fd_sc_hd__nand2_1 _5981_ (.A(_2559_),
    .B(_2557_),
    .Y(_2560_));
 sky130_fd_sc_hd__nor2_1 _5982_ (.A(_2499_),
    .B(_2492_),
    .Y(_2561_));
 sky130_fd_sc_hd__nand2_1 _5983_ (.A(_2476_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2562_));
 sky130_fd_sc_hd__o21ai_1 _5984_ (.A1(_2441_),
    .A2(_2476_),
    .B1(_2562_),
    .Y(_2563_));
 sky130_fd_sc_hd__nand3_1 _5985_ (.A(_2561_),
    .B(_2563_),
    .C(_2533_),
    .Y(_2564_));
 sky130_fd_sc_hd__nand3_1 _5986_ (.A(_2478_),
    .B(_2533_),
    .C(_2495_),
    .Y(_2565_));
 sky130_fd_sc_hd__nand2_1 _5987_ (.A(_2476_),
    .B(_2428_),
    .Y(_2566_));
 sky130_fd_sc_hd__o21ai_1 _5988_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .A2(_2476_),
    .B1(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__nand2_1 _5989_ (.A(_2565_),
    .B(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__nand3_1 _5990_ (.A(_2564_),
    .B(_2568_),
    .C(_2479_),
    .Y(_2569_));
 sky130_fd_sc_hd__nand2_1 _5991_ (.A(_2540_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2570_));
 sky130_fd_sc_hd__or2_1 _5992_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(_2540_),
    .X(_2571_));
 sky130_fd_sc_hd__and3_1 _5993_ (.A(_2502_),
    .B(_2570_),
    .C(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__or2_1 _5994_ (.A(_2421_),
    .B(_2427_),
    .X(_2573_));
 sky130_fd_sc_hd__nor2_1 _5995_ (.A(_2426_),
    .B(_2514_),
    .Y(_2574_));
 sky130_fd_sc_hd__inv_2 _5996_ (.A(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__nand2_1 _5997_ (.A(_2573_),
    .B(_2575_),
    .Y(_2576_));
 sky130_fd_sc_hd__mux2_1 _5998_ (.A0(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .A1(_2506_),
    .S(_2513_),
    .X(_2577_));
 sky130_fd_sc_hd__a22o_1 _5999_ (.A1(_2457_),
    .A2(_2576_),
    .B1(_2550_),
    .B2(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__nor2_1 _6000_ (.A(_2572_),
    .B(_2578_),
    .Y(_2579_));
 sky130_fd_sc_hd__a21oi_1 _6001_ (.A1(_2569_),
    .A2(_2579_),
    .B1(_2485_),
    .Y(_2580_));
 sky130_fd_sc_hd__nand2_1 _6002_ (.A(_2560_),
    .B(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__nand2_1 _6003_ (.A(_2569_),
    .B(_2579_),
    .Y(_2582_));
 sky130_fd_sc_hd__nand2_1 _6004_ (.A(_2582_),
    .B(_2749_),
    .Y(_2583_));
 sky130_fd_sc_hd__nand3_1 _6005_ (.A(_2559_),
    .B(_2557_),
    .C(_2583_),
    .Y(_2584_));
 sky130_fd_sc_hd__nand2_1 _6006_ (.A(_2581_),
    .B(_2584_),
    .Y(_2585_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(_2585_),
    .B(_2525_),
    .Y(_2586_));
 sky130_fd_sc_hd__or2_1 _6008_ (.A(_2529_),
    .B(_2555_),
    .X(_2587_));
 sky130_fd_sc_hd__nand2_1 _6009_ (.A(net20),
    .B(net21),
    .Y(_2588_));
 sky130_fd_sc_hd__a21oi_1 _6010_ (.A1(_2586_),
    .A2(_2587_),
    .B1(_2588_),
    .Y(_2589_));
 sky130_fd_sc_hd__nand3_1 _6011_ (.A(_2586_),
    .B(_2588_),
    .C(_2587_),
    .Y(_2590_));
 sky130_fd_sc_hd__nand2_1 _6012_ (.A(_2590_),
    .B(_2407_),
    .Y(_2591_));
 sky130_fd_sc_hd__nor2_1 _6013_ (.A(_2589_),
    .B(_2591_),
    .Y(\egd_top.exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__or3_1 _6014_ (.A(_2485_),
    .B(_2410_),
    .C(_2433_),
    .X(_2592_));
 sky130_fd_sc_hd__inv_2 _6015_ (.A(_2592_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__or3_1 _6016_ (.A(_2485_),
    .B(_2410_),
    .C(_2454_),
    .X(_2593_));
 sky130_fd_sc_hd__inv_2 _6017_ (.A(_2593_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__or3_1 _6018_ (.A(_2485_),
    .B(_2410_),
    .C(_2462_),
    .X(_2594_));
 sky130_fd_sc_hd__inv_2 _6019_ (.A(_2594_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__nor2_1 _6020_ (.A(\egd_top.BitStream_buffer.pc_reg[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2595_));
 sky130_fd_sc_hd__nand2_1 _6021_ (.A(\egd_top.BitStream_buffer.pc_reg[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2596_));
 sky130_fd_sc_hd__and2b_1 _6022_ (.A_N(_2595_),
    .B(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__or2_1 _6023_ (.A(\egd_top.BitStream_buffer.pc_reg[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .X(_2598_));
 sky130_fd_sc_hd__nand2_1 _6024_ (.A(\egd_top.BitStream_buffer.pc_reg[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2599_));
 sky130_fd_sc_hd__nand2_2 _6025_ (.A(_2598_),
    .B(_2599_),
    .Y(_2600_));
 sky130_fd_sc_hd__o21ai_4 _6026_ (.A1(_2750_),
    .A2(_2600_),
    .B1(_2599_),
    .Y(_2601_));
 sky130_fd_sc_hd__or2_1 _6027_ (.A(\egd_top.BitStream_buffer.pc_reg[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .X(_2602_));
 sky130_fd_sc_hd__nand2_1 _6028_ (.A(\egd_top.BitStream_buffer.pc_reg[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2603_));
 sky130_fd_sc_hd__a21bo_1 _6029_ (.A1(_2601_),
    .A2(_2602_),
    .B1_N(_2603_),
    .X(_2604_));
 sky130_fd_sc_hd__xor2_2 _6030_ (.A(_2597_),
    .B(_2604_),
    .X(\egd_top.BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__and2_2 _6031_ (.A(_2602_),
    .B(_2603_),
    .X(_2605_));
 sky130_fd_sc_hd__xor2_4 _6032_ (.A(_2605_),
    .B(_2601_),
    .X(\egd_top.BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__o21ai_1 _6033_ (.A1(\egd_top.BitStream_buffer.pc_reg[3] ),
    .A2(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .B1(_2604_),
    .Y(_2606_));
 sky130_fd_sc_hd__nand2_1 _6034_ (.A(_2606_),
    .B(_2596_),
    .Y(_2607_));
 sky130_fd_sc_hd__or2_1 _6035_ (.A(\egd_top.BitStream_buffer.pc_reg[4] ),
    .B(_2607_),
    .X(_2608_));
 sky130_fd_sc_hd__nand2_1 _6036_ (.A(_2607_),
    .B(\egd_top.BitStream_buffer.pc_reg[4] ),
    .Y(_2609_));
 sky130_fd_sc_hd__and2_1 _6037_ (.A(_2608_),
    .B(_2609_),
    .X(_2610_));
 sky130_fd_sc_hd__clkbuf_2 _6038_ (.A(_2610_),
    .X(\egd_top.BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__xor2_4 _6039_ (.A(_2750_),
    .B(_2600_),
    .X(\egd_top.BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__inv_2 _6040_ (.A(\egd_top.BitStream_buffer.pc_reg[5] ),
    .Y(_2611_));
 sky130_fd_sc_hd__or2_2 _6041_ (.A(_2611_),
    .B(_2609_),
    .X(_2612_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_2609_),
    .B(_2611_),
    .Y(_2613_));
 sky130_fd_sc_hd__and2_1 _6043_ (.A(_2612_),
    .B(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__clkbuf_2 _6044_ (.A(_2614_),
    .X(\egd_top.BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__xnor2_4 _6045_ (.A(\egd_top.BitStream_buffer.pc_reg[6] ),
    .B(_2612_),
    .Y(\egd_top.BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nand2_1 _6046_ (.A(_2586_),
    .B(_2587_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_1 _6047_ (.A(_2567_),
    .B(_2533_),
    .Y(_2615_));
 sky130_fd_sc_hd__nand2_1 _6048_ (.A(_2476_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2616_));
 sky130_fd_sc_hd__o21ai_2 _6049_ (.A1(_2443_),
    .A2(_2476_),
    .B1(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__inv_2 _6050_ (.A(_2617_),
    .Y(_2618_));
 sky130_fd_sc_hd__o21ai_1 _6051_ (.A1(_2530_),
    .A2(_2615_),
    .B1(_2618_),
    .Y(_2619_));
 sky130_fd_sc_hd__nor2_1 _6052_ (.A(_2530_),
    .B(_2615_),
    .Y(_2620_));
 sky130_fd_sc_hd__nand2_1 _6053_ (.A(_2620_),
    .B(_2617_),
    .Y(_2621_));
 sky130_fd_sc_hd__nand3_1 _6054_ (.A(_2619_),
    .B(_2621_),
    .C(_2479_),
    .Y(_2622_));
 sky130_fd_sc_hd__nor2_1 _6055_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2574_),
    .Y(_2623_));
 sky130_fd_sc_hd__nor2_1 _6056_ (.A(_2420_),
    .B(_2575_),
    .Y(_2624_));
 sky130_fd_sc_hd__nand2_1 _6057_ (.A(_2513_),
    .B(_2503_),
    .Y(_2625_));
 sky130_fd_sc_hd__xor2_1 _6058_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__o32a_1 _6059_ (.A1(_2623_),
    .A2(_2624_),
    .A3(_2458_),
    .B1(_2463_),
    .B2(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__nand2_2 _6060_ (.A(_2622_),
    .B(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__nand2_2 _6061_ (.A(_2628_),
    .B(_2749_),
    .Y(_2629_));
 sky130_fd_sc_hd__nor2_1 _6062_ (.A(_2557_),
    .B(_2580_),
    .Y(_2630_));
 sky130_fd_sc_hd__nor2_1 _6063_ (.A(_2629_),
    .B(_2630_),
    .Y(_2631_));
 sky130_fd_sc_hd__nand2_1 _6064_ (.A(_2629_),
    .B(_2583_),
    .Y(_2632_));
 sky130_fd_sc_hd__nor2_1 _6065_ (.A(_2557_),
    .B(_2632_),
    .Y(_2633_));
 sky130_fd_sc_hd__o21a_1 _6066_ (.A1(_2631_),
    .A2(_2633_),
    .B1(_2482_),
    .X(_2634_));
 sky130_fd_sc_hd__nor2_1 _6067_ (.A(_2524_),
    .B(_2555_),
    .Y(_2635_));
 sky130_fd_sc_hd__nand2_1 _6068_ (.A(_2580_),
    .B(_2635_),
    .Y(_2636_));
 sky130_fd_sc_hd__nor2_1 _6069_ (.A(_2629_),
    .B(_2636_),
    .Y(_2637_));
 sky130_fd_sc_hd__and2_1 _6070_ (.A(_2636_),
    .B(_2629_),
    .X(_2638_));
 sky130_fd_sc_hd__o21ai_1 _6071_ (.A1(_2637_),
    .A2(_2638_),
    .B1(_2483_),
    .Y(_2639_));
 sky130_fd_sc_hd__nand2_1 _6072_ (.A(_2639_),
    .B(_2525_),
    .Y(_2640_));
 sky130_fd_sc_hd__inv_2 _6073_ (.A(_2529_),
    .Y(_2641_));
 sky130_fd_sc_hd__nand2_1 _6074_ (.A(_2582_),
    .B(_2641_),
    .Y(_2642_));
 sky130_fd_sc_hd__o21ai_2 _6075_ (.A1(_2634_),
    .A2(_2640_),
    .B1(_2642_),
    .Y(net23));
 sky130_fd_sc_hd__nand2_1 _6076_ (.A(_2633_),
    .B(_2482_),
    .Y(_2643_));
 sky130_fd_sc_hd__o21ai_1 _6077_ (.A1(_2629_),
    .A2(_2636_),
    .B1(_2483_),
    .Y(_2644_));
 sky130_fd_sc_hd__nand2_1 _6078_ (.A(_2643_),
    .B(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__nor2_1 _6079_ (.A(_2537_),
    .B(_2563_),
    .Y(_2646_));
 sky130_fd_sc_hd__nand3_1 _6080_ (.A(_2646_),
    .B(_2561_),
    .C(_2618_),
    .Y(_2647_));
 sky130_fd_sc_hd__a21oi_2 _6081_ (.A1(_2476_),
    .A2(_2441_),
    .B1(_2421_),
    .Y(_2648_));
 sky130_fd_sc_hd__inv_2 _6082_ (.A(_2648_),
    .Y(_2649_));
 sky130_fd_sc_hd__nand2_1 _6083_ (.A(_2647_),
    .B(_2649_),
    .Y(_2650_));
 sky130_fd_sc_hd__nand3_1 _6084_ (.A(_2620_),
    .B(_2648_),
    .C(_2618_),
    .Y(_2651_));
 sky130_fd_sc_hd__nand3_1 _6085_ (.A(_2650_),
    .B(_2651_),
    .C(_2479_),
    .Y(_2652_));
 sky130_fd_sc_hd__nor2_1 _6086_ (.A(_2506_),
    .B(_2575_),
    .Y(_2653_));
 sky130_fd_sc_hd__a211o_1 _6087_ (.A1(_2417_),
    .A2(_2575_),
    .B1(_2653_),
    .C1(_2458_),
    .X(_2654_));
 sky130_fd_sc_hd__nand2_1 _6088_ (.A(_2652_),
    .B(_2654_),
    .Y(_2655_));
 sky130_fd_sc_hd__nand2_1 _6089_ (.A(_2655_),
    .B(_2749_),
    .Y(_2656_));
 sky130_fd_sc_hd__nand2_1 _6090_ (.A(_2645_),
    .B(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__inv_2 _6091_ (.A(_2656_),
    .Y(_2658_));
 sky130_fd_sc_hd__nand3_1 _6092_ (.A(_2643_),
    .B(_2644_),
    .C(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__nand3_1 _6093_ (.A(_2657_),
    .B(_2659_),
    .C(_2525_),
    .Y(_2660_));
 sky130_fd_sc_hd__nand2_1 _6094_ (.A(_2628_),
    .B(_2641_),
    .Y(_2661_));
 sky130_fd_sc_hd__nand2_1 _6095_ (.A(_2660_),
    .B(_2661_),
    .Y(net24));
 sky130_fd_sc_hd__nand3_1 _6096_ (.A(_2655_),
    .B(_2749_),
    .C(_2628_),
    .Y(_2662_));
 sky130_fd_sc_hd__inv_2 _6097_ (.A(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__nor3_1 _6098_ (.A(_2555_),
    .B(_2524_),
    .C(_2583_),
    .Y(_2664_));
 sky130_fd_sc_hd__nand2_1 _6099_ (.A(_2663_),
    .B(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__nor2_1 _6100_ (.A(_2648_),
    .B(_2617_),
    .Y(_2666_));
 sky130_fd_sc_hd__nand2_1 _6101_ (.A(_2620_),
    .B(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__o21ai_2 _6102_ (.A1(_2443_),
    .A2(_2489_),
    .B1(_2420_),
    .Y(_2668_));
 sky130_fd_sc_hd__inv_2 _6103_ (.A(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__nand2_1 _6104_ (.A(_2667_),
    .B(_2669_),
    .Y(_2670_));
 sky130_fd_sc_hd__nand3_1 _6105_ (.A(_2620_),
    .B(_2666_),
    .C(_2668_),
    .Y(_2671_));
 sky130_fd_sc_hd__nand3_1 _6106_ (.A(_2670_),
    .B(_2479_),
    .C(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__nor2_2 _6107_ (.A(_2485_),
    .B(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__inv_2 _6108_ (.A(_2673_),
    .Y(_2674_));
 sky130_fd_sc_hd__nand2_1 _6109_ (.A(_2665_),
    .B(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__nand3_1 _6110_ (.A(_2663_),
    .B(_2664_),
    .C(_2673_),
    .Y(_2676_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_2675_),
    .B(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__nand2_1 _6112_ (.A(_2677_),
    .B(_2483_),
    .Y(_2678_));
 sky130_fd_sc_hd__nand3_1 _6113_ (.A(_2630_),
    .B(_2629_),
    .C(_2656_),
    .Y(_2679_));
 sky130_fd_sc_hd__nand2_1 _6114_ (.A(_2679_),
    .B(_2673_),
    .Y(_2680_));
 sky130_fd_sc_hd__a21oi_1 _6115_ (.A1(_2655_),
    .A2(_2749_),
    .B1(_2673_),
    .Y(_2681_));
 sky130_fd_sc_hd__nand2_1 _6116_ (.A(_2633_),
    .B(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__nand2_1 _6117_ (.A(_2680_),
    .B(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__nand2_1 _6118_ (.A(_2683_),
    .B(_2482_),
    .Y(_2684_));
 sky130_fd_sc_hd__nand3_1 _6119_ (.A(_2678_),
    .B(_2684_),
    .C(_2525_),
    .Y(_2685_));
 sky130_fd_sc_hd__nand2_1 _6120_ (.A(_2655_),
    .B(_2641_),
    .Y(_2686_));
 sky130_fd_sc_hd__nand2_1 _6121_ (.A(_2685_),
    .B(_2686_),
    .Y(net25));
 sky130_fd_sc_hd__nand3_1 _6122_ (.A(_2637_),
    .B(_2673_),
    .C(_2658_),
    .Y(_2687_));
 sky130_fd_sc_hd__or2_1 _6123_ (.A(_2668_),
    .B(_2667_),
    .X(_2688_));
 sky130_fd_sc_hd__nand2_1 _6124_ (.A(_2688_),
    .B(_2476_),
    .Y(_2689_));
 sky130_fd_sc_hd__inv_2 _6125_ (.A(_2689_),
    .Y(_2690_));
 sky130_fd_sc_hd__nand2_1 _6126_ (.A(_2690_),
    .B(_2749_),
    .Y(_2691_));
 sky130_fd_sc_hd__nand2_1 _6127_ (.A(_2687_),
    .B(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__nand2_1 _6128_ (.A(_2692_),
    .B(_2483_),
    .Y(_2693_));
 sky130_fd_sc_hd__inv_2 _6129_ (.A(_2691_),
    .Y(_2694_));
 sky130_fd_sc_hd__nand2_1 _6130_ (.A(_2682_),
    .B(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__nor2_1 _6131_ (.A(_2486_),
    .B(_2481_),
    .Y(_2696_));
 sky130_fd_sc_hd__nand2_1 _6132_ (.A(_2695_),
    .B(_2696_),
    .Y(_2697_));
 sky130_fd_sc_hd__nand2_1 _6133_ (.A(_2693_),
    .B(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__nand2_1 _6134_ (.A(_2698_),
    .B(_2525_),
    .Y(_2699_));
 sky130_fd_sc_hd__a211o_1 _6135_ (.A1(net18),
    .A2(_2410_),
    .B1(_2745_),
    .C1(_2672_),
    .X(_2700_));
 sky130_fd_sc_hd__nand2_1 _6136_ (.A(_2699_),
    .B(_2700_),
    .Y(net26));
 sky130_fd_sc_hd__a211o_1 _6137_ (.A1(net18),
    .A2(_2410_),
    .B1(_2745_),
    .C1(_2689_),
    .X(_2701_));
 sky130_fd_sc_hd__a21bo_1 _6138_ (.A1(_2525_),
    .A2(_2696_),
    .B1_N(_2701_),
    .X(net27));
 sky130_fd_sc_hd__buf_8 _6139_ (.A(net19),
    .X(_2702_));
 sky130_fd_sc_hd__inv_2 _6140_ (.A(_2702_),
    .Y(_0000_));
 sky130_fd_sc_hd__buf_4 _6141_ (.A(net19),
    .X(_2703_));
 sky130_fd_sc_hd__clkbuf_8 _6142_ (.A(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__inv_2 _6143_ (.A(_2704_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _6144_ (.A(_2704_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _6145_ (.A(_2704_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _6146_ (.A(_2704_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _6147_ (.A(_2704_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _6148_ (.A(_2704_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _6149_ (.A(_2704_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _6150_ (.A(_2704_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _6151_ (.A(_2704_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _6152_ (.A(_2704_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _6153_ (.A(_2704_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _6154_ (.A(_2704_),
    .Y(_0012_));
 sky130_fd_sc_hd__clkbuf_8 _6155_ (.A(_2703_),
    .X(_2705_));
 sky130_fd_sc_hd__inv_2 _6156_ (.A(_2705_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _6157_ (.A(_2705_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _6158_ (.A(_2705_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_1 _6159_ (.A(\egd_top.BitStream_buffer.pc[0] ),
    .B(_0000_),
    .Y(_2706_));
 sky130_fd_sc_hd__inv_2 _6160_ (.A(_2706_),
    .Y(_0177_));
 sky130_fd_sc_hd__nor2_1 _6161_ (.A(_2703_),
    .B(_2819_),
    .Y(_0178_));
 sky130_fd_sc_hd__nor2_1 _6162_ (.A(_2703_),
    .B(_2818_),
    .Y(_0179_));
 sky130_fd_sc_hd__nor2_1 _6163_ (.A(_2703_),
    .B(_2872_),
    .Y(_0180_));
 sky130_fd_sc_hd__nor2_1 _6164_ (.A(_2703_),
    .B(_2933_),
    .Y(_0181_));
 sky130_fd_sc_hd__nor2_1 _6165_ (.A(_2703_),
    .B(_2822_),
    .Y(_0182_));
 sky130_fd_sc_hd__nor2_1 _6166_ (.A(_2703_),
    .B(_2754_),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _6167_ (.A(_2705_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _6168_ (.A(_2705_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _6169_ (.A(_2705_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _6170_ (.A(_2705_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _6171_ (.A(_2705_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _6172_ (.A(_2705_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _6173_ (.A(_2705_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _6174_ (.A(_2705_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _6175_ (.A(_2705_),
    .Y(_0024_));
 sky130_fd_sc_hd__clkbuf_8 _6176_ (.A(_2702_),
    .X(_2707_));
 sky130_fd_sc_hd__inv_2 _6177_ (.A(_2707_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _6178_ (.A(_2707_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _6179_ (.A(_2707_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _6180_ (.A(_2707_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _6181_ (.A(_2707_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _6182_ (.A(_2707_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _6183_ (.A(_2707_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _6184_ (.A(_2707_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _6185_ (.A(_2707_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _6186_ (.A(_2707_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _6187_ (.A(_2707_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _6188_ (.A(_2707_),
    .Y(_0036_));
 sky130_fd_sc_hd__clkbuf_8 _6189_ (.A(_2702_),
    .X(_2708_));
 sky130_fd_sc_hd__inv_2 _6190_ (.A(_2708_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _6191_ (.A(_2708_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _6192_ (.A(_2708_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _6193_ (.A(_2708_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _6194_ (.A(_2708_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _6195_ (.A(_2708_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _6196_ (.A(_2708_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _6197_ (.A(_2708_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _6198_ (.A(_2708_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _6199_ (.A(_2708_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _6200_ (.A(_2708_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _6201_ (.A(_2708_),
    .Y(_0048_));
 sky130_fd_sc_hd__clkbuf_8 _6202_ (.A(_2702_),
    .X(_2709_));
 sky130_fd_sc_hd__inv_2 _6203_ (.A(_2709_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _6204_ (.A(_2709_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _6205_ (.A(_2709_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _6206_ (.A(_2709_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _6207_ (.A(_2709_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _6208_ (.A(_2709_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _6209_ (.A(_2709_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _6210_ (.A(_2709_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _6211_ (.A(_2709_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _6212_ (.A(_2709_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _6213_ (.A(_2709_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _6214_ (.A(_2709_),
    .Y(_0060_));
 sky130_fd_sc_hd__clkbuf_8 _6215_ (.A(_2702_),
    .X(_2710_));
 sky130_fd_sc_hd__inv_2 _6216_ (.A(_2710_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _6217_ (.A(_2710_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _6218_ (.A(_2710_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _6219_ (.A(_2710_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _6220_ (.A(_2710_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _6221_ (.A(_2710_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _6222_ (.A(_2710_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _6223_ (.A(_2710_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _6224_ (.A(_2710_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _6225_ (.A(_2710_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _6226_ (.A(_2710_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _6227_ (.A(_2710_),
    .Y(_0072_));
 sky130_fd_sc_hd__clkbuf_8 _6228_ (.A(_2702_),
    .X(_2711_));
 sky130_fd_sc_hd__inv_2 _6229_ (.A(_2711_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _6230_ (.A(_2711_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _6231_ (.A(_2711_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _6232_ (.A(_2711_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _6233_ (.A(_2711_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _6234_ (.A(_2711_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _6235_ (.A(_2711_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _6236_ (.A(_2711_),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _6237_ (.A(_2711_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _6238_ (.A(_2711_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _6239_ (.A(_2711_),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _6240_ (.A(_2711_),
    .Y(_0084_));
 sky130_fd_sc_hd__clkbuf_8 _6241_ (.A(_2702_),
    .X(_2712_));
 sky130_fd_sc_hd__inv_2 _6242_ (.A(_2712_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _6243_ (.A(_2712_),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _6244_ (.A(_2712_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _6245_ (.A(_2712_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _6246_ (.A(_2712_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _6247_ (.A(_2712_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _6248_ (.A(_2712_),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _6249_ (.A(_2712_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _6250_ (.A(_2712_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _6251_ (.A(_2712_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _6252_ (.A(_2712_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _6253_ (.A(_2712_),
    .Y(_0096_));
 sky130_fd_sc_hd__clkbuf_8 _6254_ (.A(_2702_),
    .X(_2713_));
 sky130_fd_sc_hd__inv_2 _6255_ (.A(_2713_),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _6256_ (.A(_2713_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _6257_ (.A(_2713_),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _6258_ (.A(_2713_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _6259_ (.A(_2713_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _6260_ (.A(_2713_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _6261_ (.A(_2713_),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _6262_ (.A(_2713_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _6263_ (.A(_2713_),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _6264_ (.A(_2713_),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _6265_ (.A(_2713_),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _6266_ (.A(_2713_),
    .Y(_0108_));
 sky130_fd_sc_hd__clkbuf_8 _6267_ (.A(_2702_),
    .X(_2714_));
 sky130_fd_sc_hd__inv_2 _6268_ (.A(_2714_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _6269_ (.A(_2714_),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _6270_ (.A(_2714_),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _6271_ (.A(_2714_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _6272_ (.A(_2714_),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _6273_ (.A(_2714_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _6274_ (.A(_2714_),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _6275_ (.A(_2714_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _6276_ (.A(_2714_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _6277_ (.A(_2714_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _6278_ (.A(_2714_),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _6279_ (.A(_2714_),
    .Y(_0120_));
 sky130_fd_sc_hd__clkbuf_8 _6280_ (.A(_2702_),
    .X(_2715_));
 sky130_fd_sc_hd__inv_2 _6281_ (.A(_2715_),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _6282_ (.A(_2715_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _6283_ (.A(_2715_),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _6284_ (.A(_2715_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _6285_ (.A(_2715_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _6286_ (.A(_2715_),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _6287_ (.A(_2715_),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _6288_ (.A(_2715_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _6289_ (.A(_2715_),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _6290_ (.A(_2715_),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _6291_ (.A(_2715_),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _6292_ (.A(_2715_),
    .Y(_0132_));
 sky130_fd_sc_hd__clkbuf_8 _6293_ (.A(_2702_),
    .X(_2716_));
 sky130_fd_sc_hd__inv_2 _6294_ (.A(_2716_),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _6295_ (.A(_2716_),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _6296_ (.A(_2716_),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _6297_ (.A(_2716_),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _6298_ (.A(_2716_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _6299_ (.A(_2716_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _6300_ (.A(_2716_),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _6301_ (.A(_2716_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _6302_ (.A(_2716_),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _6303_ (.A(_2716_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _6304_ (.A(_2716_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _6305_ (.A(_2716_),
    .Y(_0144_));
 sky130_fd_sc_hd__clkbuf_8 _6306_ (.A(_2702_),
    .X(_2717_));
 sky130_fd_sc_hd__inv_2 _6307_ (.A(_2717_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _6308_ (.A(_2717_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _6309_ (.A(_2717_),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _6310_ (.A(_2717_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _6311_ (.A(_2717_),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _6312_ (.A(_2717_),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _6313_ (.A(_2717_),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _6314_ (.A(_2717_),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _6315_ (.A(_2717_),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _6316_ (.A(_2717_),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _6317_ (.A(_2717_),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _6318_ (.A(_2717_),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _6319_ (.A(_2703_),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _6320_ (.A(_2703_),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _6321_ (.A(_2703_),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _6322_ (.A(_2703_),
    .Y(_0160_));
 sky130_fd_sc_hd__dfrtp_4 _6323_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0161_),
    .RESET_B(_0000_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfrtp_2 _6324_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0162_),
    .RESET_B(_0001_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfrtp_2 _6325_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0163_),
    .RESET_B(_0002_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfrtp_2 _6326_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0164_),
    .RESET_B(_0003_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfrtp_4 _6327_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0165_),
    .RESET_B(_0004_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfrtp_4 _6328_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0166_),
    .RESET_B(_0005_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfrtp_2 _6329_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0167_),
    .RESET_B(_0006_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfrtp_2 _6330_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0168_),
    .RESET_B(_0007_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfrtp_2 _6331_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0169_),
    .RESET_B(_0008_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfrtp_2 _6332_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0170_),
    .RESET_B(_0009_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfrtp_4 _6333_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0171_),
    .RESET_B(_0010_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfrtp_4 _6334_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0172_),
    .RESET_B(_0011_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfrtp_4 _6335_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0173_),
    .RESET_B(_0012_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfrtp_4 _6336_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0174_),
    .RESET_B(_0013_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfrtp_4 _6337_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0175_),
    .RESET_B(_0014_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfrtp_4 _6338_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0176_),
    .RESET_B(_0015_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_1 _6339_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0177_),
    .Q(\egd_top.BitStream_buffer.pc_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6340_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0178_),
    .Q(\egd_top.BitStream_buffer.pc_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6341_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0179_),
    .Q(\egd_top.BitStream_buffer.pc_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6342_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0180_),
    .Q(\egd_top.BitStream_buffer.pc_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6343_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0181_),
    .Q(\egd_top.BitStream_buffer.pc_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6344_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0182_),
    .Q(\egd_top.BitStream_buffer.pc_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6345_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0183_),
    .Q(\egd_top.BitStream_buffer.pc_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6346_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0184_),
    .RESET_B(_0016_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfrtp_1 _6347_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0185_),
    .RESET_B(_0017_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfrtp_1 _6348_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0186_),
    .RESET_B(_0018_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfrtp_2 _6349_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0187_),
    .RESET_B(_0019_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfrtp_1 _6350_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0188_),
    .RESET_B(_0020_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfrtp_1 _6351_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0189_),
    .RESET_B(_0021_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfrtp_1 _6352_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0190_),
    .RESET_B(_0022_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfrtp_1 _6353_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0191_),
    .RESET_B(_0023_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfrtp_2 _6354_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0192_),
    .RESET_B(_0024_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfrtp_1 _6355_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_0193_),
    .RESET_B(_0025_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfrtp_4 _6356_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0194_),
    .RESET_B(_0026_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfrtp_1 _6357_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0195_),
    .RESET_B(_0027_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfrtp_1 _6358_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0196_),
    .RESET_B(_0028_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfrtp_1 _6359_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0197_),
    .RESET_B(_0029_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfrtp_2 _6360_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0198_),
    .RESET_B(_0030_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfrtp_2 _6361_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0199_),
    .RESET_B(_0031_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfrtp_2 _6362_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0200_),
    .RESET_B(_0032_),
    .Q(\egd_top.BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6363_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0201_),
    .RESET_B(_0033_),
    .Q(\egd_top.BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6364_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_0202_),
    .RESET_B(_0034_),
    .Q(\egd_top.BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6365_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0203_),
    .RESET_B(_0035_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfrtp_4 _6366_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_0204_),
    .RESET_B(_0036_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfrtp_4 _6367_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0205_),
    .RESET_B(_0037_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfrtp_4 _6368_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0206_),
    .RESET_B(_0038_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfrtp_4 _6369_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0207_),
    .RESET_B(_0039_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfrtp_4 _6370_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0208_),
    .RESET_B(_0040_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfrtp_4 _6371_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0209_),
    .RESET_B(_0041_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfrtp_2 _6372_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_0210_),
    .RESET_B(_0042_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfrtp_2 _6373_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0211_),
    .RESET_B(_0043_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfrtp_2 _6374_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0212_),
    .RESET_B(_0044_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfrtp_2 _6375_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0213_),
    .RESET_B(_0045_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfrtp_4 _6376_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0214_),
    .RESET_B(_0046_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfrtp_2 _6377_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0215_),
    .RESET_B(_0047_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfrtp_1 _6378_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0216_),
    .RESET_B(_0048_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfrtp_1 _6379_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0217_),
    .RESET_B(_0049_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfrtp_1 _6380_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0218_),
    .RESET_B(_0050_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfrtp_1 _6381_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0219_),
    .RESET_B(_0051_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfrtp_1 _6382_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0220_),
    .RESET_B(_0052_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfrtp_1 _6383_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0221_),
    .RESET_B(_0053_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfrtp_1 _6384_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0222_),
    .RESET_B(_0054_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfrtp_1 _6385_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0223_),
    .RESET_B(_0055_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfrtp_1 _6386_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0224_),
    .RESET_B(_0056_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfrtp_4 _6387_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0225_),
    .RESET_B(_0057_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfrtp_4 _6388_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0226_),
    .RESET_B(_0058_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfrtp_4 _6389_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0227_),
    .RESET_B(_0059_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfrtp_4 _6390_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_0228_),
    .RESET_B(_0060_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfrtp_4 _6391_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0229_),
    .RESET_B(_0061_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfrtp_1 _6392_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0230_),
    .RESET_B(_0062_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfrtp_1 _6393_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0231_),
    .RESET_B(_0063_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfrtp_1 _6394_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0232_),
    .RESET_B(_0064_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfrtp_1 _6395_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0233_),
    .RESET_B(_0065_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfrtp_1 _6396_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0234_),
    .RESET_B(_0066_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfrtp_1 _6397_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0235_),
    .RESET_B(_0067_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfrtp_1 _6398_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0236_),
    .RESET_B(_0068_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfrtp_1 _6399_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_0237_),
    .RESET_B(_0069_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfrtp_1 _6400_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0238_),
    .RESET_B(_0070_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfrtp_1 _6401_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0239_),
    .RESET_B(_0071_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfrtp_1 _6402_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_0240_),
    .RESET_B(_0072_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfrtp_1 _6403_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0241_),
    .RESET_B(_0073_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfrtp_2 _6404_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0242_),
    .RESET_B(_0074_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfrtp_2 _6405_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0243_),
    .RESET_B(_0075_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfrtp_1 _6406_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0244_),
    .RESET_B(_0076_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfrtp_4 _6407_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0245_),
    .RESET_B(_0077_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfrtp_1 _6408_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0246_),
    .RESET_B(_0078_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfrtp_1 _6409_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0247_),
    .RESET_B(_0079_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfrtp_1 _6410_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0248_),
    .RESET_B(_0080_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfrtp_1 _6411_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0249_),
    .RESET_B(_0081_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfrtp_1 _6412_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0250_),
    .RESET_B(_0082_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfrtp_1 _6413_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_0251_),
    .RESET_B(_0083_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6414_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_0252_),
    .RESET_B(_0084_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfrtp_1 _6415_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0253_),
    .RESET_B(_0085_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfrtp_1 _6416_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0254_),
    .RESET_B(_0086_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfrtp_1 _6417_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0255_),
    .RESET_B(_0087_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfrtp_1 _6418_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0256_),
    .RESET_B(_0088_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfrtp_1 _6419_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0257_),
    .RESET_B(_0089_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfrtp_1 _6420_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0258_),
    .RESET_B(_0090_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfrtp_1 _6421_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0259_),
    .RESET_B(_0091_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6422_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0260_),
    .RESET_B(_0092_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6423_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0261_),
    .RESET_B(_0093_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6424_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0262_),
    .RESET_B(_0094_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6425_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0263_),
    .RESET_B(_0095_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6426_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0264_),
    .RESET_B(_0096_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6427_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0265_),
    .RESET_B(_0097_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6428_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0266_),
    .RESET_B(_0098_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfrtp_1 _6429_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0267_),
    .RESET_B(_0099_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6430_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0268_),
    .RESET_B(_0100_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6431_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0269_),
    .RESET_B(_0101_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6432_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0270_),
    .RESET_B(_0102_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6433_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0271_),
    .RESET_B(_0103_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6434_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0272_),
    .RESET_B(_0104_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6435_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0273_),
    .RESET_B(_0105_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6436_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0274_),
    .RESET_B(_0106_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6437_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0275_),
    .RESET_B(_0107_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6438_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0276_),
    .RESET_B(_0108_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6439_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0277_),
    .RESET_B(_0109_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6440_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0278_),
    .RESET_B(_0110_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6441_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0279_),
    .RESET_B(_0111_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6442_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0280_),
    .RESET_B(_0112_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6443_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0281_),
    .RESET_B(_0113_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6444_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0282_),
    .RESET_B(_0114_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6445_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0283_),
    .RESET_B(_0115_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6446_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0284_),
    .RESET_B(_0116_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6447_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0285_),
    .RESET_B(_0117_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6448_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0286_),
    .RESET_B(_0118_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6449_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0287_),
    .RESET_B(_0119_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6450_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0288_),
    .RESET_B(_0120_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6451_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0289_),
    .RESET_B(_0121_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6452_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0290_),
    .RESET_B(_0122_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6453_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0291_),
    .RESET_B(_0123_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6454_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0292_),
    .RESET_B(_0124_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6455_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0293_),
    .RESET_B(_0125_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6456_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0294_),
    .RESET_B(_0126_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6457_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0295_),
    .RESET_B(_0127_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6458_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0296_),
    .RESET_B(_0128_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6459_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0297_),
    .RESET_B(_0129_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6460_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_0298_),
    .RESET_B(_0130_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfrtp_4 _6461_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0299_),
    .RESET_B(_0131_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfrtp_4 _6462_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0300_),
    .RESET_B(_0132_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfrtp_4 _6463_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0301_),
    .RESET_B(_0133_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfrtp_2 _6464_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0302_),
    .RESET_B(_0134_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfrtp_1 _6465_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0303_),
    .RESET_B(_0135_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfrtp_1 _6466_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0304_),
    .RESET_B(_0136_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfrtp_1 _6467_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_0305_),
    .RESET_B(_0137_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfrtp_1 _6468_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0306_),
    .RESET_B(_0138_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfrtp_1 _6469_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0307_),
    .RESET_B(_0139_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfrtp_1 _6470_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0308_),
    .RESET_B(_0140_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfrtp_1 _6471_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_0309_),
    .RESET_B(_0141_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfrtp_1 _6472_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0310_),
    .RESET_B(_0142_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfrtp_1 _6473_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0311_),
    .RESET_B(_0143_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfrtp_1 _6474_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_0312_),
    .RESET_B(_0144_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfrtp_1 _6475_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0313_),
    .RESET_B(_0145_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfstp_1 _6476_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_0314_),
    .SET_B(_0146_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 _6477_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0315_),
    .RESET_B(_0147_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_4 _6478_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0316_),
    .RESET_B(_0148_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_4 _6479_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_0317_),
    .RESET_B(_0149_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _6480_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(\egd_top.BitStream_buffer.pc[0] ),
    .RESET_B(_0150_),
    .Q(\egd_top.BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6481_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(\egd_top.BitStream_buffer.pc[1] ),
    .RESET_B(_0151_),
    .Q(\egd_top.BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6482_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(\egd_top.BitStream_buffer.pc[2] ),
    .RESET_B(_0152_),
    .Q(\egd_top.BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6483_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(\egd_top.BitStream_buffer.pc[3] ),
    .RESET_B(_0153_),
    .Q(\egd_top.BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6484_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(\egd_top.BitStream_buffer.pc[4] ),
    .RESET_B(_0154_),
    .Q(\egd_top.BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6485_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(\egd_top.BitStream_buffer.pc[5] ),
    .RESET_B(_0155_),
    .Q(\egd_top.BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6486_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(\egd_top.BitStream_buffer.pc[6] ),
    .RESET_B(_0156_),
    .Q(\egd_top.BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6487_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0318_),
    .RESET_B(_0157_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_4 _6488_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0319_),
    .RESET_B(_0158_),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_2 _6489_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0320_),
    .RESET_B(_0159_),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_2 _6490_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_0321_),
    .RESET_B(_0160_),
    .Q(net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__buf_4 input1 (.A(la_data_in_47_32[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(la_data_in_47_32[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(la_data_in_47_32[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(la_data_in_47_32[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(la_data_in_47_32[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(la_data_in_47_32[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 input15 (.A(la_data_in_47_32[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(la_data_in_47_32[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(la_data_in_49_48[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(la_data_in_49_48[1]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(wb_rst_i),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(la_data_in_47_32[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_8 input3 (.A(la_data_in_47_32[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(la_data_in_47_32[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(la_data_in_47_32[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(la_data_in_47_32[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(la_data_in_47_32[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(la_data_in_47_32[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(la_data_in_47_32[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 max_cap35 (.A(_2900_),
    .X(net35));
 sky130_fd_sc_hd__buf_4 max_cap36 (.A(_2834_),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 max_cap38 (.A(_2821_),
    .X(net38));
 sky130_fd_sc_hd__buf_4 max_cap39 (.A(\egd_top.BitStream_buffer.pc[3] ),
    .X(net39));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(la_data_out_15_8[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(la_data_out_15_8[1]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(la_data_out_15_8[2]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(la_data_out_15_8[3]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(la_data_out_15_8[4]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(la_data_out_15_8[5]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(la_data_out_15_8[6]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_data_out_15_8[7]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(la_data_out_18_16[0]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(la_data_out_18_16[1]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(la_data_out_18_16[2]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(la_data_out_22_19[0]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(la_data_out_22_19[1]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(la_data_out_22_19[2]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(la_data_out_22_19[3]));
 sky130_fd_sc_hd__buf_2 wire37 (.A(_2829_),
    .X(net37));
endmodule

