// This is the unpowered netlist.
module egd_top_wrapper (la_data_in_64,
    la_data_in_65,
    la_oenb_64,
    wb_clk_i,
    la_data_in_47_32,
    la_data_in_49_48,
    la_data_out_15_8,
    la_data_out_18_16,
    la_data_out_22_19);
 input la_data_in_64;
 input la_data_in_65;
 input la_oenb_64;
 input wb_clk_i;
 input [15:0] la_data_in_47_32;
 input [1:0] la_data_in_49_48;
 output [7:0] la_data_out_15_8;
 output [2:0] la_data_out_18_16;
 output [3:0] la_data_out_22_19;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire clknet_0__2956_;
 wire clknet_0__2957_;
 wire clknet_0__2958_;
 wire clknet_0__2961_;
 wire clknet_0__2964_;
 wire clknet_0__2967_;
 wire clknet_0__2970_;
 wire clknet_0__2973_;
 wire clknet_0__2976_;
 wire clknet_0__2979_;
 wire clknet_0__2982_;
 wire clknet_0__2985_;
 wire clknet_0__2988_;
 wire clknet_0__2991_;
 wire clknet_0__2994_;
 wire clknet_0__2997_;
 wire clknet_0__3000_;
 wire clknet_0__3003_;
 wire clknet_1_0__leaf__2956_;
 wire clknet_1_0__leaf__2957_;
 wire clknet_1_0__leaf__2958_;
 wire clknet_1_0__leaf__2961_;
 wire clknet_1_0__leaf__2964_;
 wire clknet_1_0__leaf__2967_;
 wire clknet_1_0__leaf__2970_;
 wire clknet_1_0__leaf__2973_;
 wire clknet_1_0__leaf__2976_;
 wire clknet_1_0__leaf__2979_;
 wire clknet_1_0__leaf__2982_;
 wire clknet_1_0__leaf__2985_;
 wire clknet_1_0__leaf__2988_;
 wire clknet_1_0__leaf__2991_;
 wire clknet_1_0__leaf__2994_;
 wire clknet_1_0__leaf__2997_;
 wire clknet_1_0__leaf__3000_;
 wire clknet_1_0__leaf__3003_;
 wire clknet_1_1__leaf__2956_;
 wire clknet_1_1__leaf__2957_;
 wire clknet_1_1__leaf__2958_;
 wire clknet_1_1__leaf__2961_;
 wire clknet_1_1__leaf__2964_;
 wire clknet_1_1__leaf__2967_;
 wire clknet_1_1__leaf__2970_;
 wire clknet_1_1__leaf__2973_;
 wire clknet_1_1__leaf__2976_;
 wire clknet_1_1__leaf__2979_;
 wire clknet_1_1__leaf__2982_;
 wire clknet_1_1__leaf__2985_;
 wire clknet_1_1__leaf__2988_;
 wire clknet_1_1__leaf__2991_;
 wire clknet_1_1__leaf__2994_;
 wire clknet_1_1__leaf__2997_;
 wire clknet_1_1__leaf__3000_;
 wire clknet_1_1__leaf__3003_;
 wire \egd_top.BitStream_buffer.BS_buffer[0] ;
 wire \egd_top.BitStream_buffer.BS_buffer[100] ;
 wire \egd_top.BitStream_buffer.BS_buffer[101] ;
 wire \egd_top.BitStream_buffer.BS_buffer[102] ;
 wire \egd_top.BitStream_buffer.BS_buffer[103] ;
 wire \egd_top.BitStream_buffer.BS_buffer[104] ;
 wire \egd_top.BitStream_buffer.BS_buffer[105] ;
 wire \egd_top.BitStream_buffer.BS_buffer[106] ;
 wire \egd_top.BitStream_buffer.BS_buffer[107] ;
 wire \egd_top.BitStream_buffer.BS_buffer[108] ;
 wire \egd_top.BitStream_buffer.BS_buffer[109] ;
 wire \egd_top.BitStream_buffer.BS_buffer[10] ;
 wire \egd_top.BitStream_buffer.BS_buffer[110] ;
 wire \egd_top.BitStream_buffer.BS_buffer[111] ;
 wire \egd_top.BitStream_buffer.BS_buffer[112] ;
 wire \egd_top.BitStream_buffer.BS_buffer[113] ;
 wire \egd_top.BitStream_buffer.BS_buffer[114] ;
 wire \egd_top.BitStream_buffer.BS_buffer[115] ;
 wire \egd_top.BitStream_buffer.BS_buffer[116] ;
 wire \egd_top.BitStream_buffer.BS_buffer[117] ;
 wire \egd_top.BitStream_buffer.BS_buffer[118] ;
 wire \egd_top.BitStream_buffer.BS_buffer[119] ;
 wire \egd_top.BitStream_buffer.BS_buffer[11] ;
 wire \egd_top.BitStream_buffer.BS_buffer[120] ;
 wire \egd_top.BitStream_buffer.BS_buffer[121] ;
 wire \egd_top.BitStream_buffer.BS_buffer[122] ;
 wire \egd_top.BitStream_buffer.BS_buffer[123] ;
 wire \egd_top.BitStream_buffer.BS_buffer[124] ;
 wire \egd_top.BitStream_buffer.BS_buffer[125] ;
 wire \egd_top.BitStream_buffer.BS_buffer[126] ;
 wire \egd_top.BitStream_buffer.BS_buffer[127] ;
 wire \egd_top.BitStream_buffer.BS_buffer[12] ;
 wire \egd_top.BitStream_buffer.BS_buffer[13] ;
 wire \egd_top.BitStream_buffer.BS_buffer[14] ;
 wire \egd_top.BitStream_buffer.BS_buffer[15] ;
 wire \egd_top.BitStream_buffer.BS_buffer[16] ;
 wire \egd_top.BitStream_buffer.BS_buffer[17] ;
 wire \egd_top.BitStream_buffer.BS_buffer[18] ;
 wire \egd_top.BitStream_buffer.BS_buffer[19] ;
 wire \egd_top.BitStream_buffer.BS_buffer[1] ;
 wire \egd_top.BitStream_buffer.BS_buffer[20] ;
 wire \egd_top.BitStream_buffer.BS_buffer[21] ;
 wire \egd_top.BitStream_buffer.BS_buffer[22] ;
 wire \egd_top.BitStream_buffer.BS_buffer[23] ;
 wire \egd_top.BitStream_buffer.BS_buffer[24] ;
 wire \egd_top.BitStream_buffer.BS_buffer[25] ;
 wire \egd_top.BitStream_buffer.BS_buffer[26] ;
 wire \egd_top.BitStream_buffer.BS_buffer[27] ;
 wire \egd_top.BitStream_buffer.BS_buffer[28] ;
 wire \egd_top.BitStream_buffer.BS_buffer[29] ;
 wire \egd_top.BitStream_buffer.BS_buffer[2] ;
 wire \egd_top.BitStream_buffer.BS_buffer[30] ;
 wire \egd_top.BitStream_buffer.BS_buffer[31] ;
 wire \egd_top.BitStream_buffer.BS_buffer[32] ;
 wire \egd_top.BitStream_buffer.BS_buffer[33] ;
 wire \egd_top.BitStream_buffer.BS_buffer[34] ;
 wire \egd_top.BitStream_buffer.BS_buffer[35] ;
 wire \egd_top.BitStream_buffer.BS_buffer[36] ;
 wire \egd_top.BitStream_buffer.BS_buffer[37] ;
 wire \egd_top.BitStream_buffer.BS_buffer[38] ;
 wire \egd_top.BitStream_buffer.BS_buffer[39] ;
 wire \egd_top.BitStream_buffer.BS_buffer[3] ;
 wire \egd_top.BitStream_buffer.BS_buffer[40] ;
 wire \egd_top.BitStream_buffer.BS_buffer[41] ;
 wire \egd_top.BitStream_buffer.BS_buffer[42] ;
 wire \egd_top.BitStream_buffer.BS_buffer[43] ;
 wire \egd_top.BitStream_buffer.BS_buffer[44] ;
 wire \egd_top.BitStream_buffer.BS_buffer[45] ;
 wire \egd_top.BitStream_buffer.BS_buffer[46] ;
 wire \egd_top.BitStream_buffer.BS_buffer[47] ;
 wire \egd_top.BitStream_buffer.BS_buffer[48] ;
 wire \egd_top.BitStream_buffer.BS_buffer[49] ;
 wire \egd_top.BitStream_buffer.BS_buffer[4] ;
 wire \egd_top.BitStream_buffer.BS_buffer[50] ;
 wire \egd_top.BitStream_buffer.BS_buffer[51] ;
 wire \egd_top.BitStream_buffer.BS_buffer[52] ;
 wire \egd_top.BitStream_buffer.BS_buffer[53] ;
 wire \egd_top.BitStream_buffer.BS_buffer[54] ;
 wire \egd_top.BitStream_buffer.BS_buffer[55] ;
 wire \egd_top.BitStream_buffer.BS_buffer[56] ;
 wire \egd_top.BitStream_buffer.BS_buffer[57] ;
 wire \egd_top.BitStream_buffer.BS_buffer[58] ;
 wire \egd_top.BitStream_buffer.BS_buffer[59] ;
 wire \egd_top.BitStream_buffer.BS_buffer[5] ;
 wire \egd_top.BitStream_buffer.BS_buffer[60] ;
 wire \egd_top.BitStream_buffer.BS_buffer[61] ;
 wire \egd_top.BitStream_buffer.BS_buffer[62] ;
 wire \egd_top.BitStream_buffer.BS_buffer[63] ;
 wire \egd_top.BitStream_buffer.BS_buffer[64] ;
 wire \egd_top.BitStream_buffer.BS_buffer[65] ;
 wire \egd_top.BitStream_buffer.BS_buffer[66] ;
 wire \egd_top.BitStream_buffer.BS_buffer[67] ;
 wire \egd_top.BitStream_buffer.BS_buffer[68] ;
 wire \egd_top.BitStream_buffer.BS_buffer[69] ;
 wire \egd_top.BitStream_buffer.BS_buffer[6] ;
 wire \egd_top.BitStream_buffer.BS_buffer[70] ;
 wire \egd_top.BitStream_buffer.BS_buffer[71] ;
 wire \egd_top.BitStream_buffer.BS_buffer[72] ;
 wire \egd_top.BitStream_buffer.BS_buffer[73] ;
 wire \egd_top.BitStream_buffer.BS_buffer[74] ;
 wire \egd_top.BitStream_buffer.BS_buffer[75] ;
 wire \egd_top.BitStream_buffer.BS_buffer[76] ;
 wire \egd_top.BitStream_buffer.BS_buffer[77] ;
 wire \egd_top.BitStream_buffer.BS_buffer[78] ;
 wire \egd_top.BitStream_buffer.BS_buffer[79] ;
 wire \egd_top.BitStream_buffer.BS_buffer[7] ;
 wire \egd_top.BitStream_buffer.BS_buffer[80] ;
 wire \egd_top.BitStream_buffer.BS_buffer[81] ;
 wire \egd_top.BitStream_buffer.BS_buffer[82] ;
 wire \egd_top.BitStream_buffer.BS_buffer[83] ;
 wire \egd_top.BitStream_buffer.BS_buffer[84] ;
 wire \egd_top.BitStream_buffer.BS_buffer[85] ;
 wire \egd_top.BitStream_buffer.BS_buffer[86] ;
 wire \egd_top.BitStream_buffer.BS_buffer[87] ;
 wire \egd_top.BitStream_buffer.BS_buffer[88] ;
 wire \egd_top.BitStream_buffer.BS_buffer[89] ;
 wire \egd_top.BitStream_buffer.BS_buffer[8] ;
 wire \egd_top.BitStream_buffer.BS_buffer[90] ;
 wire \egd_top.BitStream_buffer.BS_buffer[91] ;
 wire \egd_top.BitStream_buffer.BS_buffer[92] ;
 wire \egd_top.BitStream_buffer.BS_buffer[93] ;
 wire \egd_top.BitStream_buffer.BS_buffer[94] ;
 wire \egd_top.BitStream_buffer.BS_buffer[95] ;
 wire \egd_top.BitStream_buffer.BS_buffer[96] ;
 wire \egd_top.BitStream_buffer.BS_buffer[97] ;
 wire \egd_top.BitStream_buffer.BS_buffer[98] ;
 wire \egd_top.BitStream_buffer.BS_buffer[99] ;
 wire \egd_top.BitStream_buffer.BS_buffer[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[10] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[11] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[12] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[13] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[14] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[15] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[1] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[2] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[3] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[4] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[5] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[6] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[7] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[8] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_valid_n ;
 wire \egd_top.BitStream_buffer.buffer_index[4] ;
 wire \egd_top.BitStream_buffer.buffer_index[5] ;
 wire \egd_top.BitStream_buffer.buffer_index[6] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[1] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[2] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[3] ;
 wire \egd_top.BitStream_buffer.pc[1] ;
 wire \egd_top.BitStream_buffer.pc[2] ;
 wire \egd_top.BitStream_buffer.pc[3] ;
 wire \egd_top.BitStream_buffer.pc[4] ;
 wire \egd_top.BitStream_buffer.pc[5] ;
 wire \egd_top.BitStream_buffer.pc[6] ;
 wire \egd_top.BitStream_buffer.pc_previous[0] ;
 wire \egd_top.BitStream_buffer.pc_previous[1] ;
 wire \egd_top.BitStream_buffer.pc_previous[2] ;
 wire \egd_top.BitStream_buffer.pc_previous[3] ;
 wire \egd_top.BitStream_buffer.pc_previous[4] ;
 wire \egd_top.BitStream_buffer.pc_previous[5] ;
 wire \egd_top.BitStream_buffer.pc_previous[6] ;
 wire \egd_top.exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1794_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_2032_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net4));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3444_ (.A(net35),
    .Y(_3004_));
 sky130_fd_sc_hd__nand2_1 _3445_ (.A(net34),
    .B(net33),
    .Y(_3005_));
 sky130_fd_sc_hd__inv_2 _3446_ (.A(net36),
    .Y(_3006_));
 sky130_fd_sc_hd__o21ai_1 _3447_ (.A1(_3004_),
    .A2(_3005_),
    .B1(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__clkbuf_4 _3448_ (.A(net20),
    .X(_3008_));
 sky130_fd_sc_hd__buf_2 _3449_ (.A(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__and2_1 _3450_ (.A(_3007_),
    .B(_3009_),
    .X(_3010_));
 sky130_fd_sc_hd__clkbuf_1 _3451_ (.A(_3010_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_1 _3452_ (.A1(_3004_),
    .A2(_3005_),
    .B1(_3007_),
    .X(_3011_));
 sky130_fd_sc_hd__nand2_1 _3453_ (.A(net36),
    .B(net35),
    .Y(_3012_));
 sky130_fd_sc_hd__inv_2 _3454_ (.A(net20),
    .Y(_3013_));
 sky130_fd_sc_hd__a21oi_1 _3455_ (.A1(_3011_),
    .A2(_3012_),
    .B1(_3013_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _3456_ (.A(net33),
    .Y(_3014_));
 sky130_fd_sc_hd__nor2_1 _3457_ (.A(net35),
    .B(net34),
    .Y(_3015_));
 sky130_fd_sc_hd__nor2_1 _3458_ (.A(_3006_),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__nor2_1 _3459_ (.A(_3014_),
    .B(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__a21o_1 _3460_ (.A1(_3017_),
    .A2(net34),
    .B1(_3013_),
    .X(_3018_));
 sky130_fd_sc_hd__o21ba_1 _3461_ (.A1(net34),
    .A2(_3017_),
    .B1_N(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__clkbuf_1 _3462_ (.A(_3019_),
    .X(_0319_));
 sky130_fd_sc_hd__inv_2 _3463_ (.A(_3016_),
    .Y(_3020_));
 sky130_fd_sc_hd__nor2_1 _3464_ (.A(net33),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__or3_1 _3465_ (.A(_3013_),
    .B(_3017_),
    .C(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__inv_2 _3466_ (.A(_3022_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _3467_ (.A(net32),
    .Y(_3023_));
 sky130_fd_sc_hd__nor2_1 _3468_ (.A(net31),
    .B(net30),
    .Y(_3024_));
 sky130_fd_sc_hd__nor2_1 _3469_ (.A(_3023_),
    .B(_3024_),
    .Y(_3025_));
 sky130_fd_sc_hd__a21o_1 _3470_ (.A1(net31),
    .A2(net30),
    .B1(net32),
    .X(_3026_));
 sky130_fd_sc_hd__and2b_1 _3471_ (.A_N(_3025_),
    .B(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__inv_2 _3472_ (.A(net31),
    .Y(_3028_));
 sky130_fd_sc_hd__nand2_4 _3473_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3029_));
 sky130_fd_sc_hd__inv_2 _3474_ (.A(net18),
    .Y(_3030_));
 sky130_fd_sc_hd__inv_2 _3475_ (.A(net17),
    .Y(_3031_));
 sky130_fd_sc_hd__nand2_4 _3476_ (.A(_3030_),
    .B(_3031_),
    .Y(_3032_));
 sky130_fd_sc_hd__or2_1 _3477_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__nand2_4 _3478_ (.A(_3032_),
    .B(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_3034_));
 sky130_fd_sc_hd__nand2_2 _3479_ (.A(_3033_),
    .B(_3034_),
    .Y(_3035_));
 sky130_fd_sc_hd__inv_2 _3480_ (.A(_3035_),
    .Y(_3036_));
 sky130_fd_sc_hd__nand2_2 _3481_ (.A(_3036_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3037_));
 sky130_fd_sc_hd__nor2_4 _3482_ (.A(_3029_),
    .B(_3037_),
    .Y(_3038_));
 sky130_fd_sc_hd__inv_2 _3483_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_3039_));
 sky130_fd_sc_hd__and3_1 _3484_ (.A(_3039_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3040_));
 sky130_fd_sc_hd__and2_2 _3485_ (.A(_3038_),
    .B(_3040_),
    .X(_3041_));
 sky130_fd_sc_hd__nor2_1 _3486_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__inv_2 _3487_ (.A(_3024_),
    .Y(_3043_));
 sky130_fd_sc_hd__nor2_1 _3488_ (.A(net32),
    .B(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__inv_2 _3489_ (.A(net39),
    .Y(_3045_));
 sky130_fd_sc_hd__inv_2 _3490_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_3046_));
 sky130_fd_sc_hd__and3_1 _3491_ (.A(_3045_),
    .B(_3046_),
    .C(net37),
    .X(_3047_));
 sky130_fd_sc_hd__nand3_1 _3492_ (.A(_3042_),
    .B(_3044_),
    .C(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__nor2_1 _3493_ (.A(_3025_),
    .B(_3044_),
    .Y(_3049_));
 sky130_fd_sc_hd__inv_2 _3494_ (.A(_3049_),
    .Y(_3050_));
 sky130_fd_sc_hd__nand2_1 _3495_ (.A(_3048_),
    .B(_3050_),
    .Y(_3051_));
 sky130_fd_sc_hd__inv_2 _3496_ (.A(net37),
    .Y(_3052_));
 sky130_fd_sc_hd__and3_1 _3497_ (.A(_3052_),
    .B(_3045_),
    .C(_3046_),
    .X(_3053_));
 sky130_fd_sc_hd__and2b_1 _3498_ (.A_N(_3053_),
    .B(\egd_top.BitStream_buffer.pc_previous[6] ),
    .X(_3054_));
 sky130_fd_sc_hd__and4_1 _3499_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(\egd_top.BitStream_buffer.pc_previous[1] ),
    .C(\egd_top.BitStream_buffer.pc_previous[2] ),
    .D(\egd_top.BitStream_buffer.pc_previous[3] ),
    .X(_3055_));
 sky130_fd_sc_hd__a31o_1 _3500_ (.A1(_3055_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .A3(\egd_top.BitStream_buffer.pc_previous[5] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[6] ),
    .X(_3056_));
 sky130_fd_sc_hd__nand2_1 _3501_ (.A(_3042_),
    .B(_3056_),
    .Y(_3057_));
 sky130_fd_sc_hd__o21ai_1 _3502_ (.A1(_3039_),
    .A2(_3054_),
    .B1(_3057_),
    .Y(_3058_));
 sky130_fd_sc_hd__and2_1 _3503_ (.A(_3058_),
    .B(_3044_),
    .X(_3059_));
 sky130_fd_sc_hd__a311o_1 _3504_ (.A1(net32),
    .A2(_3028_),
    .A3(net30),
    .B1(_3051_),
    .C1(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__and4_1 _3505_ (.A(_3004_),
    .B(_3014_),
    .C(net36),
    .D(net34),
    .X(_3061_));
 sky130_fd_sc_hd__nand2_2 _3506_ (.A(_3060_),
    .B(_3061_),
    .Y(_3062_));
 sky130_fd_sc_hd__clkbuf_4 _3507_ (.A(_3008_),
    .X(_3063_));
 sky130_fd_sc_hd__nand2_1 _3508_ (.A(_3062_),
    .B(_3023_),
    .Y(_3064_));
 sky130_fd_sc_hd__o211a_1 _3509_ (.A1(_3027_),
    .A2(_3062_),
    .B1(_3063_),
    .C1(_3064_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _3510_ (.A(_3024_),
    .B(_3026_),
    .Y(_3065_));
 sky130_fd_sc_hd__nand2_1 _3511_ (.A(_3062_),
    .B(_3028_),
    .Y(_3066_));
 sky130_fd_sc_hd__o211a_1 _3512_ (.A1(_3065_),
    .A2(_3062_),
    .B1(_3063_),
    .C1(_3066_),
    .X(_0316_));
 sky130_fd_sc_hd__o21ai_1 _3513_ (.A1(net30),
    .A2(_3050_),
    .B1(_3048_),
    .Y(_3067_));
 sky130_fd_sc_hd__o21bai_1 _3514_ (.A1(_3059_),
    .A2(_3067_),
    .B1_N(_3062_),
    .Y(_3068_));
 sky130_fd_sc_hd__nand2_1 _3515_ (.A(_3062_),
    .B(net30),
    .Y(_3069_));
 sky130_fd_sc_hd__a21oi_1 _3516_ (.A1(_3068_),
    .A2(_3069_),
    .B1(_3013_),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _3517_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .Y(_3070_));
 sky130_fd_sc_hd__clkbuf_4 _3518_ (.A(_3070_),
    .X(_3071_));
 sky130_fd_sc_hd__o21ai_1 _3519_ (.A1(_3071_),
    .A2(_3061_),
    .B1(_3063_),
    .Y(_0314_));
 sky130_fd_sc_hd__clkbuf_4 _3520_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .X(_3072_));
 sky130_fd_sc_hd__nand2_1 _3521_ (.A(_3023_),
    .B(_3028_),
    .Y(_3073_));
 sky130_fd_sc_hd__nand2_1 _3522_ (.A(net32),
    .B(net31),
    .Y(_3074_));
 sky130_fd_sc_hd__nand2_1 _3523_ (.A(_3015_),
    .B(_3006_),
    .Y(_3075_));
 sky130_fd_sc_hd__a22o_4 _3524_ (.A1(_3073_),
    .A2(_3074_),
    .B1(_3020_),
    .B2(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__nand2_1 _3525_ (.A(_3076_),
    .B(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_3077_));
 sky130_fd_sc_hd__or2_1 _3526_ (.A(_3045_),
    .B(_3077_),
    .X(_3078_));
 sky130_fd_sc_hd__or2_1 _3527_ (.A(_3052_),
    .B(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__clkbuf_4 _3528_ (.A(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__clkbuf_4 _3529_ (.A(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(net7),
    .A1(_3072_),
    .S(_3081_),
    .X(_3082_));
 sky130_fd_sc_hd__and2_1 _3531_ (.A(_3082_),
    .B(_3009_),
    .X(_3083_));
 sky130_fd_sc_hd__clkbuf_1 _3532_ (.A(_3083_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_4 _3533_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_3084_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(net6),
    .A1(_3084_),
    .S(_3081_),
    .X(_3085_));
 sky130_fd_sc_hd__and2_1 _3535_ (.A(_3085_),
    .B(_3009_),
    .X(_3086_));
 sky130_fd_sc_hd__clkbuf_1 _3536_ (.A(_3086_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_4 _3537_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .X(_3087_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(net5),
    .A1(_3087_),
    .S(_3081_),
    .X(_3088_));
 sky130_fd_sc_hd__and2_1 _3539_ (.A(_3088_),
    .B(_3009_),
    .X(_3089_));
 sky130_fd_sc_hd__clkbuf_1 _3540_ (.A(_3089_),
    .X(_0311_));
 sky130_fd_sc_hd__buf_2 _3541_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .X(_3090_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(net4),
    .A1(_3090_),
    .S(_3081_),
    .X(_3091_));
 sky130_fd_sc_hd__and2_1 _3543_ (.A(_3091_),
    .B(_3009_),
    .X(_3092_));
 sky130_fd_sc_hd__clkbuf_1 _3544_ (.A(_3092_),
    .X(_0310_));
 sky130_fd_sc_hd__buf_2 _3545_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .X(_3093_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(net3),
    .A1(_3093_),
    .S(_3081_),
    .X(_3094_));
 sky130_fd_sc_hd__buf_4 _3547_ (.A(net20),
    .X(_3095_));
 sky130_fd_sc_hd__clkbuf_2 _3548_ (.A(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__and2_1 _3549_ (.A(_3094_),
    .B(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__clkbuf_1 _3550_ (.A(_3097_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_2 _3551_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .X(_3098_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(net2),
    .A1(_3098_),
    .S(_3081_),
    .X(_3099_));
 sky130_fd_sc_hd__and2_1 _3553_ (.A(_3099_),
    .B(_3096_),
    .X(_3100_));
 sky130_fd_sc_hd__clkbuf_1 _3554_ (.A(_3100_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_2 _3555_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .X(_3101_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(net16),
    .A1(_3101_),
    .S(_3081_),
    .X(_3102_));
 sky130_fd_sc_hd__and2_1 _3557_ (.A(_3102_),
    .B(_3096_),
    .X(_3103_));
 sky130_fd_sc_hd__clkbuf_1 _3558_ (.A(_3103_),
    .X(_0307_));
 sky130_fd_sc_hd__buf_2 _3559_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_3104_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(net15),
    .A1(_3104_),
    .S(_3081_),
    .X(_3105_));
 sky130_fd_sc_hd__and2_1 _3561_ (.A(_3105_),
    .B(_3096_),
    .X(_3106_));
 sky130_fd_sc_hd__clkbuf_1 _3562_ (.A(_3106_),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_4 _3563_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_3107_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(net14),
    .A1(_3107_),
    .S(_3081_),
    .X(_3108_));
 sky130_fd_sc_hd__and2_1 _3565_ (.A(_3108_),
    .B(_3096_),
    .X(_3109_));
 sky130_fd_sc_hd__clkbuf_1 _3566_ (.A(_3109_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_2 _3567_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_3110_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(net13),
    .A1(_3110_),
    .S(_3080_),
    .X(_3111_));
 sky130_fd_sc_hd__and2_1 _3569_ (.A(_3111_),
    .B(_3096_),
    .X(_3112_));
 sky130_fd_sc_hd__clkbuf_1 _3570_ (.A(_3112_),
    .X(_0304_));
 sky130_fd_sc_hd__buf_2 _3571_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_3113_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(net12),
    .A1(_3113_),
    .S(_3080_),
    .X(_3114_));
 sky130_fd_sc_hd__and2_1 _3573_ (.A(_3114_),
    .B(_3096_),
    .X(_3115_));
 sky130_fd_sc_hd__clkbuf_1 _3574_ (.A(_3115_),
    .X(_0303_));
 sky130_fd_sc_hd__buf_2 _3575_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .X(_3116_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(net11),
    .A1(_3116_),
    .S(_3080_),
    .X(_3117_));
 sky130_fd_sc_hd__and2_1 _3577_ (.A(_3117_),
    .B(_3096_),
    .X(_3118_));
 sky130_fd_sc_hd__clkbuf_1 _3578_ (.A(_3118_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_2 _3579_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_3119_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(net10),
    .A1(_3119_),
    .S(_3080_),
    .X(_3120_));
 sky130_fd_sc_hd__and2_1 _3581_ (.A(_3120_),
    .B(_3096_),
    .X(_3121_));
 sky130_fd_sc_hd__clkbuf_1 _3582_ (.A(_3121_),
    .X(_0301_));
 sky130_fd_sc_hd__buf_2 _3583_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_3122_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(net9),
    .A1(_3122_),
    .S(_3080_),
    .X(_3123_));
 sky130_fd_sc_hd__and2_1 _3585_ (.A(_3123_),
    .B(_3096_),
    .X(_3124_));
 sky130_fd_sc_hd__clkbuf_1 _3586_ (.A(_3124_),
    .X(_0300_));
 sky130_fd_sc_hd__buf_2 _3587_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_3125_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(net8),
    .A1(_3125_),
    .S(_3080_),
    .X(_3126_));
 sky130_fd_sc_hd__clkbuf_2 _3589_ (.A(_3095_),
    .X(_3127_));
 sky130_fd_sc_hd__and2_1 _3590_ (.A(_3126_),
    .B(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__clkbuf_1 _3591_ (.A(_3128_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_2 _3592_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_3129_));
 sky130_fd_sc_hd__mux2_1 _3593_ (.A0(net1),
    .A1(_3129_),
    .S(_3080_),
    .X(_3130_));
 sky130_fd_sc_hd__and2_1 _3594_ (.A(_3130_),
    .B(_3127_),
    .X(_3131_));
 sky130_fd_sc_hd__clkbuf_1 _3595_ (.A(_3131_),
    .X(_0298_));
 sky130_fd_sc_hd__buf_2 _3596_ (.A(_3008_),
    .X(_3132_));
 sky130_fd_sc_hd__o21ai_1 _3597_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_3133_));
 sky130_fd_sc_hd__buf_2 _3598_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .X(_3134_));
 sky130_fd_sc_hd__clkbuf_4 _3599_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .X(_3135_));
 sky130_fd_sc_hd__inv_2 _3600_ (.A(_3135_),
    .Y(_3136_));
 sky130_fd_sc_hd__inv_2 _3601_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3137_));
 sky130_fd_sc_hd__nand2_2 _3602_ (.A(_3035_),
    .B(_3137_),
    .Y(_3138_));
 sky130_fd_sc_hd__inv_2 _3603_ (.A(_3138_),
    .Y(_3139_));
 sky130_fd_sc_hd__inv_2 _3604_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_3140_));
 sky130_fd_sc_hd__and3_1 _3605_ (.A(_3139_),
    .B(_3140_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3141_));
 sky130_fd_sc_hd__clkbuf_4 _3606_ (.A(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__inv_2 _3607_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_3143_));
 sky130_fd_sc_hd__and3_2 _3608_ (.A(_3039_),
    .B(_3143_),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_3144_));
 sky130_fd_sc_hd__buf_2 _3609_ (.A(_3144_),
    .X(_3145_));
 sky130_fd_sc_hd__nand2_2 _3610_ (.A(_3142_),
    .B(_3145_),
    .Y(_3146_));
 sky130_fd_sc_hd__buf_2 _3611_ (.A(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__nand2_2 _3612_ (.A(_3036_),
    .B(_3137_),
    .Y(_3148_));
 sky130_fd_sc_hd__inv_2 _3613_ (.A(_3148_),
    .Y(_3149_));
 sky130_fd_sc_hd__and3_1 _3614_ (.A(_3149_),
    .B(_3140_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3150_));
 sky130_fd_sc_hd__clkbuf_4 _3615_ (.A(_3150_),
    .X(_3151_));
 sky130_fd_sc_hd__and2_1 _3616_ (.A(_3151_),
    .B(_3145_),
    .X(_3152_));
 sky130_fd_sc_hd__clkbuf_2 _3617_ (.A(_3152_),
    .X(_3153_));
 sky130_fd_sc_hd__buf_4 _3618_ (.A(_3153_),
    .X(_3154_));
 sky130_fd_sc_hd__clkbuf_4 _3619_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .X(_3155_));
 sky130_fd_sc_hd__nand2_1 _3620_ (.A(_3154_),
    .B(_3155_),
    .Y(_3156_));
 sky130_fd_sc_hd__nand2_2 _3621_ (.A(_3035_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3157_));
 sky130_fd_sc_hd__inv_2 _3622_ (.A(_3157_),
    .Y(_3158_));
 sky130_fd_sc_hd__and3_2 _3623_ (.A(_3158_),
    .B(_3140_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3159_));
 sky130_fd_sc_hd__and2_2 _3624_ (.A(_3159_),
    .B(_3144_),
    .X(_3160_));
 sky130_fd_sc_hd__buf_2 _3625_ (.A(_3160_),
    .X(_3161_));
 sky130_fd_sc_hd__inv_2 _3626_ (.A(_3037_),
    .Y(_3162_));
 sky130_fd_sc_hd__and3_1 _3627_ (.A(_3162_),
    .B(_3140_),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3163_));
 sky130_fd_sc_hd__buf_6 _3628_ (.A(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__and2_2 _3629_ (.A(_3164_),
    .B(_3144_),
    .X(_3165_));
 sky130_fd_sc_hd__buf_2 _3630_ (.A(_3165_),
    .X(_3166_));
 sky130_fd_sc_hd__clkbuf_4 _3631_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .X(_3167_));
 sky130_fd_sc_hd__a22o_1 _3632_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .B1(_3166_),
    .B2(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__inv_2 _3633_ (.A(_3168_),
    .Y(_3169_));
 sky130_fd_sc_hd__o211a_1 _3634_ (.A1(_3136_),
    .A2(_3147_),
    .B1(_3156_),
    .C1(_3169_),
    .X(_3170_));
 sky130_fd_sc_hd__inv_2 _3635_ (.A(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3171_));
 sky130_fd_sc_hd__nand2_4 _3636_ (.A(_3140_),
    .B(_3171_),
    .Y(_3172_));
 sky130_fd_sc_hd__nor2_4 _3637_ (.A(_3172_),
    .B(_3138_),
    .Y(_3173_));
 sky130_fd_sc_hd__and2_1 _3638_ (.A(_3173_),
    .B(_3145_),
    .X(_3174_));
 sky130_fd_sc_hd__clkbuf_2 _3639_ (.A(_3174_),
    .X(_3175_));
 sky130_fd_sc_hd__clkbuf_4 _3640_ (.A(_3175_),
    .X(_3176_));
 sky130_fd_sc_hd__buf_2 _3641_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .X(_3177_));
 sky130_fd_sc_hd__nor2_4 _3642_ (.A(_3172_),
    .B(_3148_),
    .Y(_3178_));
 sky130_fd_sc_hd__and2_1 _3643_ (.A(_3178_),
    .B(_3145_),
    .X(_3179_));
 sky130_fd_sc_hd__clkbuf_2 _3644_ (.A(_3179_),
    .X(_3180_));
 sky130_fd_sc_hd__clkbuf_4 _3645_ (.A(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__clkbuf_4 _3646_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .X(_3182_));
 sky130_fd_sc_hd__inv_2 _3647_ (.A(_3182_),
    .Y(_3183_));
 sky130_fd_sc_hd__nor2_4 _3648_ (.A(_3172_),
    .B(_3157_),
    .Y(_3184_));
 sky130_fd_sc_hd__nand2_2 _3649_ (.A(_3184_),
    .B(_3145_),
    .Y(_3185_));
 sky130_fd_sc_hd__clkbuf_4 _3650_ (.A(_3185_),
    .X(_3186_));
 sky130_fd_sc_hd__nor2_2 _3651_ (.A(_3172_),
    .B(_3037_),
    .Y(_3187_));
 sky130_fd_sc_hd__and2_1 _3652_ (.A(_3187_),
    .B(_3145_),
    .X(_3188_));
 sky130_fd_sc_hd__clkbuf_2 _3653_ (.A(_3188_),
    .X(_3189_));
 sky130_fd_sc_hd__buf_2 _3654_ (.A(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__clkbuf_4 _3655_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .X(_3191_));
 sky130_fd_sc_hd__nand2_1 _3656_ (.A(_3190_),
    .B(_3191_),
    .Y(_3192_));
 sky130_fd_sc_hd__o21ai_1 _3657_ (.A1(_3183_),
    .A2(_3186_),
    .B1(_3192_),
    .Y(_3193_));
 sky130_fd_sc_hd__a221oi_1 _3658_ (.A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .A2(_3176_),
    .B1(_3177_),
    .B2(_3181_),
    .C1(_3193_),
    .Y(_3194_));
 sky130_fd_sc_hd__clkbuf_4 _3659_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .X(_3195_));
 sky130_fd_sc_hd__inv_2 _3660_ (.A(_3195_),
    .Y(_3196_));
 sky130_fd_sc_hd__and3_1 _3661_ (.A(_3162_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3171_),
    .X(_3197_));
 sky130_fd_sc_hd__buf_6 _3662_ (.A(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__nand2_2 _3663_ (.A(_3198_),
    .B(_3145_),
    .Y(_3199_));
 sky130_fd_sc_hd__buf_2 _3664_ (.A(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__and3_2 _3665_ (.A(_3158_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3171_),
    .X(_3201_));
 sky130_fd_sc_hd__and2_1 _3666_ (.A(_3201_),
    .B(_3144_),
    .X(_3202_));
 sky130_fd_sc_hd__clkbuf_2 _3667_ (.A(_3202_),
    .X(_3203_));
 sky130_fd_sc_hd__buf_2 _3668_ (.A(_3203_),
    .X(_3204_));
 sky130_fd_sc_hd__clkbuf_4 _3669_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .X(_3205_));
 sky130_fd_sc_hd__nand2_1 _3670_ (.A(_3204_),
    .B(_3205_),
    .Y(_3206_));
 sky130_fd_sc_hd__and3_1 _3671_ (.A(_3139_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3171_),
    .X(_3207_));
 sky130_fd_sc_hd__buf_4 _3672_ (.A(_3207_),
    .X(_3208_));
 sky130_fd_sc_hd__and2_1 _3673_ (.A(_3208_),
    .B(_3144_),
    .X(_3209_));
 sky130_fd_sc_hd__clkbuf_2 _3674_ (.A(_3209_),
    .X(_3210_));
 sky130_fd_sc_hd__buf_2 _3675_ (.A(_3210_),
    .X(_3211_));
 sky130_fd_sc_hd__clkbuf_4 _3676_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .X(_3212_));
 sky130_fd_sc_hd__nand2_1 _3677_ (.A(_3211_),
    .B(_3212_),
    .Y(_3213_));
 sky130_fd_sc_hd__clkbuf_4 _3678_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .X(_3214_));
 sky130_fd_sc_hd__inv_2 _3679_ (.A(_3214_),
    .Y(_3215_));
 sky130_fd_sc_hd__and3_1 _3680_ (.A(_3149_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3171_),
    .X(_3216_));
 sky130_fd_sc_hd__buf_4 _3681_ (.A(_3216_),
    .X(_3217_));
 sky130_fd_sc_hd__nand2_2 _3682_ (.A(_3217_),
    .B(_3145_),
    .Y(_3218_));
 sky130_fd_sc_hd__clkbuf_2 _3683_ (.A(_3218_),
    .X(_3219_));
 sky130_fd_sc_hd__or2_1 _3684_ (.A(_3215_),
    .B(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__o2111a_1 _3685_ (.A1(_3196_),
    .A2(_3200_),
    .B1(_3206_),
    .C1(_3213_),
    .D1(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__buf_2 _3686_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_3222_));
 sky130_fd_sc_hd__nor2_2 _3687_ (.A(_3029_),
    .B(_3157_),
    .Y(_3223_));
 sky130_fd_sc_hd__and2_1 _3688_ (.A(_3223_),
    .B(_3145_),
    .X(_3224_));
 sky130_fd_sc_hd__clkbuf_2 _3689_ (.A(_3224_),
    .X(_3225_));
 sky130_fd_sc_hd__buf_2 _3690_ (.A(_3225_),
    .X(_3226_));
 sky130_fd_sc_hd__buf_2 _3691_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_3227_));
 sky130_fd_sc_hd__and2_1 _3692_ (.A(_3038_),
    .B(_3145_),
    .X(_3228_));
 sky130_fd_sc_hd__clkbuf_2 _3693_ (.A(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__buf_2 _3694_ (.A(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__nor2_4 _3695_ (.A(_3029_),
    .B(_3148_),
    .Y(_3231_));
 sky130_fd_sc_hd__and2_1 _3696_ (.A(_3231_),
    .B(_3144_),
    .X(_3232_));
 sky130_fd_sc_hd__clkbuf_2 _3697_ (.A(_3232_),
    .X(_3233_));
 sky130_fd_sc_hd__buf_2 _3698_ (.A(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__clkbuf_4 _3699_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_3235_));
 sky130_fd_sc_hd__nand2_1 _3700_ (.A(_3234_),
    .B(_3235_),
    .Y(_3236_));
 sky130_fd_sc_hd__nor2_4 _3701_ (.A(_3029_),
    .B(_3138_),
    .Y(_3237_));
 sky130_fd_sc_hd__and2_1 _3702_ (.A(_3237_),
    .B(_3144_),
    .X(_3238_));
 sky130_fd_sc_hd__clkbuf_2 _3703_ (.A(_3238_),
    .X(_3239_));
 sky130_fd_sc_hd__buf_2 _3704_ (.A(_3239_),
    .X(_3240_));
 sky130_fd_sc_hd__buf_2 _3705_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_3241_));
 sky130_fd_sc_hd__nand2_1 _3706_ (.A(_3240_),
    .B(_3241_),
    .Y(_3242_));
 sky130_fd_sc_hd__nand2_1 _3707_ (.A(_3236_),
    .B(_3242_),
    .Y(_3243_));
 sky130_fd_sc_hd__a221oi_1 _3708_ (.A1(_3222_),
    .A2(_3226_),
    .B1(_3227_),
    .B2(_3230_),
    .C1(_3243_),
    .Y(_3244_));
 sky130_fd_sc_hd__and4_1 _3709_ (.A(_3170_),
    .B(_3194_),
    .C(_3221_),
    .D(_3244_),
    .X(_3245_));
 sky130_fd_sc_hd__clkbuf_4 _3710_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_3246_));
 sky130_fd_sc_hd__inv_2 _3711_ (.A(_3246_),
    .Y(_3247_));
 sky130_fd_sc_hd__inv_2 _3712_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_3248_));
 sky130_fd_sc_hd__and3_2 _3713_ (.A(_3039_),
    .B(_3248_),
    .C(_3143_),
    .X(_3249_));
 sky130_fd_sc_hd__buf_4 _3714_ (.A(_3249_),
    .X(_3250_));
 sky130_fd_sc_hd__nand2_2 _3715_ (.A(_3217_),
    .B(_3250_),
    .Y(_3251_));
 sky130_fd_sc_hd__clkbuf_4 _3716_ (.A(_3251_),
    .X(_3252_));
 sky130_fd_sc_hd__and2_1 _3717_ (.A(_3201_),
    .B(_3249_),
    .X(_3253_));
 sky130_fd_sc_hd__clkbuf_2 _3718_ (.A(_3253_),
    .X(_3254_));
 sky130_fd_sc_hd__buf_2 _3719_ (.A(_3254_),
    .X(_3255_));
 sky130_fd_sc_hd__clkbuf_4 _3720_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_3256_));
 sky130_fd_sc_hd__nand2_1 _3721_ (.A(_3255_),
    .B(_3256_),
    .Y(_3257_));
 sky130_fd_sc_hd__and2_1 _3722_ (.A(_3208_),
    .B(_3249_),
    .X(_3258_));
 sky130_fd_sc_hd__clkbuf_2 _3723_ (.A(_3258_),
    .X(_3259_));
 sky130_fd_sc_hd__buf_2 _3724_ (.A(_3259_),
    .X(_3260_));
 sky130_fd_sc_hd__buf_2 _3725_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_3261_));
 sky130_fd_sc_hd__nand2_1 _3726_ (.A(_3260_),
    .B(_3261_),
    .Y(_3262_));
 sky130_fd_sc_hd__inv_2 _3727_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_3263_));
 sky130_fd_sc_hd__nand2_1 _3728_ (.A(_3198_),
    .B(_3250_),
    .Y(_3264_));
 sky130_fd_sc_hd__buf_2 _3729_ (.A(_3264_),
    .X(_3265_));
 sky130_fd_sc_hd__or2_1 _3730_ (.A(_3263_),
    .B(_3265_),
    .X(_3266_));
 sky130_fd_sc_hd__o2111a_1 _3731_ (.A1(_3247_),
    .A2(_3252_),
    .B1(_3257_),
    .C1(_3262_),
    .D1(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__inv_2 _3732_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_3268_));
 sky130_fd_sc_hd__nand2_2 _3733_ (.A(_3164_),
    .B(_3250_),
    .Y(_3269_));
 sky130_fd_sc_hd__clkbuf_4 _3734_ (.A(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__and2_1 _3735_ (.A(_3159_),
    .B(_3249_),
    .X(_3271_));
 sky130_fd_sc_hd__clkbuf_2 _3736_ (.A(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__clkbuf_4 _3737_ (.A(_3272_),
    .X(_3273_));
 sky130_fd_sc_hd__nand2_1 _3738_ (.A(_3273_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_3274_));
 sky130_fd_sc_hd__and2_1 _3739_ (.A(_3142_),
    .B(_3249_),
    .X(_3275_));
 sky130_fd_sc_hd__clkbuf_2 _3740_ (.A(_3275_),
    .X(_3276_));
 sky130_fd_sc_hd__buf_4 _3741_ (.A(_3276_),
    .X(_3277_));
 sky130_fd_sc_hd__nand2_1 _3742_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_3278_));
 sky130_fd_sc_hd__inv_2 _3743_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_3279_));
 sky130_fd_sc_hd__nand2_1 _3744_ (.A(_3151_),
    .B(_3250_),
    .Y(_3280_));
 sky130_fd_sc_hd__buf_2 _3745_ (.A(_3280_),
    .X(_3281_));
 sky130_fd_sc_hd__or2_1 _3746_ (.A(_3279_),
    .B(_3281_),
    .X(_3282_));
 sky130_fd_sc_hd__o2111a_1 _3747_ (.A1(_3268_),
    .A2(_3270_),
    .B1(_3274_),
    .C1(_3278_),
    .D1(_3282_),
    .X(_3283_));
 sky130_fd_sc_hd__clkbuf_4 _3748_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_3284_));
 sky130_fd_sc_hd__inv_2 _3749_ (.A(_3284_),
    .Y(_3285_));
 sky130_fd_sc_hd__nand2_2 _3750_ (.A(_3184_),
    .B(_3250_),
    .Y(_3286_));
 sky130_fd_sc_hd__buf_2 _3751_ (.A(_3286_),
    .X(_3287_));
 sky130_fd_sc_hd__inv_2 _3752_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_3288_));
 sky130_fd_sc_hd__nand2_2 _3753_ (.A(_3178_),
    .B(_3250_),
    .Y(_3289_));
 sky130_fd_sc_hd__buf_2 _3754_ (.A(_3289_),
    .X(_3290_));
 sky130_fd_sc_hd__clkbuf_4 _3755_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_3291_));
 sky130_fd_sc_hd__inv_2 _3756_ (.A(_3291_),
    .Y(_3292_));
 sky130_fd_sc_hd__nand2_1 _3757_ (.A(_3187_),
    .B(_3250_),
    .Y(_3293_));
 sky130_fd_sc_hd__clkbuf_2 _3758_ (.A(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__or2_1 _3759_ (.A(_3292_),
    .B(_3294_),
    .X(_3295_));
 sky130_fd_sc_hd__o221a_1 _3760_ (.A1(_3285_),
    .A2(_3287_),
    .B1(_3288_),
    .B2(_3290_),
    .C1(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__and2_1 _3761_ (.A(_3223_),
    .B(_3249_),
    .X(_3297_));
 sky130_fd_sc_hd__clkbuf_2 _3762_ (.A(_3297_),
    .X(_3298_));
 sky130_fd_sc_hd__buf_2 _3763_ (.A(_3298_),
    .X(_3299_));
 sky130_fd_sc_hd__and2_1 _3764_ (.A(_3038_),
    .B(_3249_),
    .X(_3300_));
 sky130_fd_sc_hd__clkbuf_2 _3765_ (.A(_3300_),
    .X(_3301_));
 sky130_fd_sc_hd__buf_2 _3766_ (.A(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__inv_2 _3767_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_3303_));
 sky130_fd_sc_hd__nand2_2 _3768_ (.A(_3237_),
    .B(_3250_),
    .Y(_3304_));
 sky130_fd_sc_hd__buf_2 _3769_ (.A(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__inv_2 _3770_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_3306_));
 sky130_fd_sc_hd__nand2_2 _3771_ (.A(_3231_),
    .B(_3250_),
    .Y(_3307_));
 sky130_fd_sc_hd__buf_2 _3772_ (.A(_3307_),
    .X(_3308_));
 sky130_fd_sc_hd__o22ai_1 _3773_ (.A1(_3303_),
    .A2(_3305_),
    .B1(_3306_),
    .B2(_3308_),
    .Y(_3309_));
 sky130_fd_sc_hd__a221oi_1 _3774_ (.A1(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .A2(_3299_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .B2(_3302_),
    .C1(_3309_),
    .Y(_3310_));
 sky130_fd_sc_hd__and4_1 _3775_ (.A(_3267_),
    .B(_3283_),
    .C(_3296_),
    .D(_3310_),
    .X(_3311_));
 sky130_fd_sc_hd__clkbuf_4 _3776_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_3312_));
 sky130_fd_sc_hd__and3_2 _3777_ (.A(_3039_),
    .B(_3248_),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3313_));
 sky130_fd_sc_hd__buf_2 _3778_ (.A(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__and2_1 _3779_ (.A(_3201_),
    .B(_3314_),
    .X(_3315_));
 sky130_fd_sc_hd__clkbuf_2 _3780_ (.A(_3315_),
    .X(_3316_));
 sky130_fd_sc_hd__buf_2 _3781_ (.A(_3316_),
    .X(_3317_));
 sky130_fd_sc_hd__clkbuf_4 _3782_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_3318_));
 sky130_fd_sc_hd__and2_1 _3783_ (.A(_3198_),
    .B(_3314_),
    .X(_3319_));
 sky130_fd_sc_hd__buf_6 _3784_ (.A(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__clkbuf_4 _3785_ (.A(_3320_),
    .X(_3321_));
 sky130_fd_sc_hd__inv_2 _3786_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_3322_));
 sky130_fd_sc_hd__nand2_2 _3787_ (.A(_3208_),
    .B(_3314_),
    .Y(_3323_));
 sky130_fd_sc_hd__buf_2 _3788_ (.A(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__clkbuf_4 _3789_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_3325_));
 sky130_fd_sc_hd__inv_2 _3790_ (.A(_3325_),
    .Y(_3326_));
 sky130_fd_sc_hd__nand2_2 _3791_ (.A(_3217_),
    .B(_3314_),
    .Y(_3327_));
 sky130_fd_sc_hd__buf_2 _3792_ (.A(_3327_),
    .X(_3328_));
 sky130_fd_sc_hd__o22ai_1 _3793_ (.A1(_3322_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3328_),
    .Y(_3329_));
 sky130_fd_sc_hd__a221oi_1 _3794_ (.A1(_3312_),
    .A2(_3317_),
    .B1(_3318_),
    .B2(_3321_),
    .C1(_3329_),
    .Y(_3330_));
 sky130_fd_sc_hd__buf_2 _3795_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_3331_));
 sky130_fd_sc_hd__and2_1 _3796_ (.A(_3159_),
    .B(_3314_),
    .X(_3332_));
 sky130_fd_sc_hd__clkbuf_2 _3797_ (.A(_3332_),
    .X(_3333_));
 sky130_fd_sc_hd__buf_4 _3798_ (.A(_3333_),
    .X(_3334_));
 sky130_fd_sc_hd__buf_2 _3799_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_3335_));
 sky130_fd_sc_hd__and2_1 _3800_ (.A(_3164_),
    .B(_3314_),
    .X(_3336_));
 sky130_fd_sc_hd__clkbuf_2 _3801_ (.A(_3336_),
    .X(_3337_));
 sky130_fd_sc_hd__buf_4 _3802_ (.A(_3337_),
    .X(_3338_));
 sky130_fd_sc_hd__and2_1 _3803_ (.A(_3151_),
    .B(_3313_),
    .X(_3339_));
 sky130_fd_sc_hd__buf_6 _3804_ (.A(_3339_),
    .X(_3340_));
 sky130_fd_sc_hd__buf_6 _3805_ (.A(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__clkbuf_4 _3806_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_3342_));
 sky130_fd_sc_hd__nand2_1 _3807_ (.A(_3341_),
    .B(_3342_),
    .Y(_3343_));
 sky130_fd_sc_hd__and2_1 _3808_ (.A(_3142_),
    .B(_3313_),
    .X(_3344_));
 sky130_fd_sc_hd__clkbuf_2 _3809_ (.A(_3344_),
    .X(_3345_));
 sky130_fd_sc_hd__buf_4 _3810_ (.A(_3345_),
    .X(_3346_));
 sky130_fd_sc_hd__clkbuf_4 _3811_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_3347_));
 sky130_fd_sc_hd__nand2_1 _3812_ (.A(_3346_),
    .B(_3347_),
    .Y(_3348_));
 sky130_fd_sc_hd__nand2_1 _3813_ (.A(_3343_),
    .B(_3348_),
    .Y(_3349_));
 sky130_fd_sc_hd__a221oi_1 _3814_ (.A1(_3331_),
    .A2(_3334_),
    .B1(_3335_),
    .B2(_3338_),
    .C1(_3349_),
    .Y(_3350_));
 sky130_fd_sc_hd__clkbuf_4 _3815_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_3351_));
 sky130_fd_sc_hd__and2_1 _3816_ (.A(_3173_),
    .B(_3313_),
    .X(_3352_));
 sky130_fd_sc_hd__clkbuf_2 _3817_ (.A(_3352_),
    .X(_3353_));
 sky130_fd_sc_hd__buf_2 _3818_ (.A(_3353_),
    .X(_3354_));
 sky130_fd_sc_hd__buf_2 _3819_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_3355_));
 sky130_fd_sc_hd__and2_1 _3820_ (.A(_3178_),
    .B(_3314_),
    .X(_3356_));
 sky130_fd_sc_hd__clkbuf_2 _3821_ (.A(_3356_),
    .X(_3357_));
 sky130_fd_sc_hd__buf_2 _3822_ (.A(_3357_),
    .X(_3358_));
 sky130_fd_sc_hd__inv_2 _3823_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_3359_));
 sky130_fd_sc_hd__nand2_2 _3824_ (.A(_3184_),
    .B(_3314_),
    .Y(_3360_));
 sky130_fd_sc_hd__clkbuf_4 _3825_ (.A(_3360_),
    .X(_3361_));
 sky130_fd_sc_hd__and2_1 _3826_ (.A(_3187_),
    .B(_3313_),
    .X(_3362_));
 sky130_fd_sc_hd__clkbuf_2 _3827_ (.A(_3362_),
    .X(_3363_));
 sky130_fd_sc_hd__buf_2 _3828_ (.A(_3363_),
    .X(_3364_));
 sky130_fd_sc_hd__clkbuf_4 _3829_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_3365_));
 sky130_fd_sc_hd__nand2_1 _3830_ (.A(_3364_),
    .B(_3365_),
    .Y(_3366_));
 sky130_fd_sc_hd__o21ai_1 _3831_ (.A1(_3359_),
    .A2(_3361_),
    .B1(_3366_),
    .Y(_3367_));
 sky130_fd_sc_hd__a221oi_1 _3832_ (.A1(_3351_),
    .A2(_3354_),
    .B1(_3355_),
    .B2(_3358_),
    .C1(_3367_),
    .Y(_3368_));
 sky130_fd_sc_hd__buf_2 _3833_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_3369_));
 sky130_fd_sc_hd__and2_1 _3834_ (.A(_3237_),
    .B(_3313_),
    .X(_3370_));
 sky130_fd_sc_hd__clkbuf_2 _3835_ (.A(_3370_),
    .X(_3371_));
 sky130_fd_sc_hd__buf_2 _3836_ (.A(_3371_),
    .X(_3372_));
 sky130_fd_sc_hd__buf_2 _3837_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_3373_));
 sky130_fd_sc_hd__and2_1 _3838_ (.A(_3231_),
    .B(_3314_),
    .X(_3374_));
 sky130_fd_sc_hd__clkbuf_2 _3839_ (.A(_3374_),
    .X(_3375_));
 sky130_fd_sc_hd__buf_2 _3840_ (.A(_3375_),
    .X(_3376_));
 sky130_fd_sc_hd__inv_2 _3841_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_3377_));
 sky130_fd_sc_hd__nand2_2 _3842_ (.A(_3038_),
    .B(_3314_),
    .Y(_3378_));
 sky130_fd_sc_hd__clkbuf_4 _3843_ (.A(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__and2_1 _3844_ (.A(_3223_),
    .B(_3313_),
    .X(_3380_));
 sky130_fd_sc_hd__clkbuf_2 _3845_ (.A(_3380_),
    .X(_3381_));
 sky130_fd_sc_hd__buf_2 _3846_ (.A(_3381_),
    .X(_3382_));
 sky130_fd_sc_hd__nand2_1 _3847_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_3383_));
 sky130_fd_sc_hd__o21ai_1 _3848_ (.A1(_3377_),
    .A2(_3379_),
    .B1(_3383_),
    .Y(_3384_));
 sky130_fd_sc_hd__a221oi_1 _3849_ (.A1(_3369_),
    .A2(_3372_),
    .B1(_3373_),
    .B2(_3376_),
    .C1(_3384_),
    .Y(_3385_));
 sky130_fd_sc_hd__and4_1 _3850_ (.A(_3330_),
    .B(_3350_),
    .C(_3368_),
    .D(_3385_),
    .X(_3386_));
 sky130_fd_sc_hd__inv_2 _3851_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_3387_));
 sky130_fd_sc_hd__buf_2 _3852_ (.A(_3040_),
    .X(_3388_));
 sky130_fd_sc_hd__nand2_2 _3853_ (.A(_3217_),
    .B(_3388_),
    .Y(_3389_));
 sky130_fd_sc_hd__buf_2 _3854_ (.A(_3389_),
    .X(_3390_));
 sky130_fd_sc_hd__and2_1 _3855_ (.A(_3201_),
    .B(_3040_),
    .X(_3391_));
 sky130_fd_sc_hd__clkbuf_2 _3856_ (.A(_3391_),
    .X(_3392_));
 sky130_fd_sc_hd__buf_2 _3857_ (.A(_3392_),
    .X(_3393_));
 sky130_fd_sc_hd__buf_2 _3858_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .X(_3394_));
 sky130_fd_sc_hd__nand2_1 _3859_ (.A(_3393_),
    .B(_3394_),
    .Y(_3395_));
 sky130_fd_sc_hd__and2_1 _3860_ (.A(_3208_),
    .B(_3388_),
    .X(_3396_));
 sky130_fd_sc_hd__clkbuf_2 _3861_ (.A(_3396_),
    .X(_3397_));
 sky130_fd_sc_hd__buf_4 _3862_ (.A(_3397_),
    .X(_3398_));
 sky130_fd_sc_hd__clkbuf_4 _3863_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_3399_));
 sky130_fd_sc_hd__nand2_1 _3864_ (.A(_3398_),
    .B(_3399_),
    .Y(_3400_));
 sky130_fd_sc_hd__inv_2 _3865_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_3401_));
 sky130_fd_sc_hd__nand2_2 _3866_ (.A(_3198_),
    .B(_3388_),
    .Y(_3402_));
 sky130_fd_sc_hd__clkbuf_2 _3867_ (.A(_3402_),
    .X(_3403_));
 sky130_fd_sc_hd__or2_1 _3868_ (.A(_3401_),
    .B(_3403_),
    .X(_3404_));
 sky130_fd_sc_hd__o2111a_1 _3869_ (.A1(_3387_),
    .A2(_3390_),
    .B1(_3395_),
    .C1(_3400_),
    .D1(_3404_),
    .X(_3405_));
 sky130_fd_sc_hd__inv_2 _3870_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .Y(_3406_));
 sky130_fd_sc_hd__nand2_2 _3871_ (.A(_3164_),
    .B(_3388_),
    .Y(_3407_));
 sky130_fd_sc_hd__clkbuf_4 _3872_ (.A(_3407_),
    .X(_3408_));
 sky130_fd_sc_hd__and2_1 _3873_ (.A(_3142_),
    .B(_3040_),
    .X(_3409_));
 sky130_fd_sc_hd__clkbuf_2 _3874_ (.A(_3409_),
    .X(_3410_));
 sky130_fd_sc_hd__buf_4 _3875_ (.A(_3410_),
    .X(_3411_));
 sky130_fd_sc_hd__nand2_1 _3876_ (.A(_3411_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_3412_));
 sky130_fd_sc_hd__and2_1 _3877_ (.A(_3159_),
    .B(_3040_),
    .X(_3413_));
 sky130_fd_sc_hd__clkbuf_2 _3878_ (.A(_3413_),
    .X(_3414_));
 sky130_fd_sc_hd__buf_2 _3879_ (.A(_3414_),
    .X(_3415_));
 sky130_fd_sc_hd__buf_2 _3880_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .X(_3416_));
 sky130_fd_sc_hd__nand2_1 _3881_ (.A(_3415_),
    .B(_3416_),
    .Y(_3417_));
 sky130_fd_sc_hd__inv_2 _3882_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_3418_));
 sky130_fd_sc_hd__nand2_1 _3883_ (.A(_3151_),
    .B(_3388_),
    .Y(_3419_));
 sky130_fd_sc_hd__clkbuf_2 _3884_ (.A(_3419_),
    .X(_3420_));
 sky130_fd_sc_hd__or2_1 _3885_ (.A(_3418_),
    .B(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__o2111a_1 _3886_ (.A1(_3406_),
    .A2(_3408_),
    .B1(_3412_),
    .C1(_3417_),
    .D1(_3421_),
    .X(_3422_));
 sky130_fd_sc_hd__buf_2 _3887_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_3423_));
 sky130_fd_sc_hd__and2_1 _3888_ (.A(_3184_),
    .B(_3388_),
    .X(_3424_));
 sky130_fd_sc_hd__clkbuf_2 _3889_ (.A(_3424_),
    .X(_3425_));
 sky130_fd_sc_hd__buf_2 _3890_ (.A(_3425_),
    .X(_3426_));
 sky130_fd_sc_hd__buf_2 _3891_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_3427_));
 sky130_fd_sc_hd__and2_1 _3892_ (.A(_3187_),
    .B(_3388_),
    .X(_3428_));
 sky130_fd_sc_hd__clkbuf_2 _3893_ (.A(_3428_),
    .X(_3429_));
 sky130_fd_sc_hd__buf_2 _3894_ (.A(_3429_),
    .X(_3430_));
 sky130_fd_sc_hd__inv_2 _3895_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .Y(_3431_));
 sky130_fd_sc_hd__nand2_2 _3896_ (.A(_3173_),
    .B(_3388_),
    .Y(_3432_));
 sky130_fd_sc_hd__clkbuf_4 _3897_ (.A(_3432_),
    .X(_3433_));
 sky130_fd_sc_hd__and2_1 _3898_ (.A(_3178_),
    .B(_3040_),
    .X(_3434_));
 sky130_fd_sc_hd__clkbuf_2 _3899_ (.A(_3434_),
    .X(_3435_));
 sky130_fd_sc_hd__buf_2 _3900_ (.A(_3435_),
    .X(_3436_));
 sky130_fd_sc_hd__nand2_1 _3901_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_3437_));
 sky130_fd_sc_hd__o21ai_1 _3902_ (.A1(_3431_),
    .A2(_3433_),
    .B1(_3437_),
    .Y(_3438_));
 sky130_fd_sc_hd__a221oi_1 _3903_ (.A1(_3423_),
    .A2(_3426_),
    .B1(_3427_),
    .B2(_3430_),
    .C1(_3438_),
    .Y(_3439_));
 sky130_fd_sc_hd__buf_2 _3904_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .X(_3440_));
 sky130_fd_sc_hd__and2_1 _3905_ (.A(_3237_),
    .B(_3388_),
    .X(_3441_));
 sky130_fd_sc_hd__clkbuf_2 _3906_ (.A(_3441_),
    .X(_3442_));
 sky130_fd_sc_hd__buf_2 _3907_ (.A(_3442_),
    .X(_3443_));
 sky130_fd_sc_hd__buf_2 _3908_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _3909_ (.A(_3231_),
    .B(_3388_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_2 _3910_ (.A(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__buf_2 _3911_ (.A(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__inv_2 _3912_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _3913_ (.A(_3041_),
    .Y(_0327_));
 sky130_fd_sc_hd__buf_2 _3914_ (.A(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__and2_1 _3915_ (.A(_3223_),
    .B(_3040_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_2 _3916_ (.A(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__buf_2 _3917_ (.A(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _3918_ (.A(_0331_),
    .B(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_0332_));
 sky130_fd_sc_hd__o21ai_1 _3919_ (.A1(_0326_),
    .A2(_0328_),
    .B1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__a221oi_1 _3920_ (.A1(_3440_),
    .A2(_3443_),
    .B1(_0322_),
    .B2(_0325_),
    .C1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__and4_1 _3921_ (.A(_3405_),
    .B(_3422_),
    .C(_3439_),
    .D(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__and4_1 _3922_ (.A(_3245_),
    .B(_3311_),
    .C(_3386_),
    .D(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_4 _3923_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_0337_));
 sky130_fd_sc_hd__and3_2 _3924_ (.A(_3248_),
    .B(_3143_),
    .C(\egd_top.BitStream_buffer.pc[6] ),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_4 _3925_ (.A(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__and2_1 _3926_ (.A(_3159_),
    .B(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_2 _3927_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_2 _3928_ (.A(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__buf_2 _3929_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_0343_));
 sky130_fd_sc_hd__and2_1 _3930_ (.A(_3164_),
    .B(_0339_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_2 _3931_ (.A(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__buf_6 _3932_ (.A(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__inv_2 _3933_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_2 _3934_ (.A(_3142_),
    .B(_0339_),
    .Y(_0348_));
 sky130_fd_sc_hd__buf_2 _3935_ (.A(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_4 _3936_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_0350_));
 sky130_fd_sc_hd__inv_2 _3937_ (.A(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_2 _3938_ (.A(_3151_),
    .B(_0339_),
    .Y(_0352_));
 sky130_fd_sc_hd__clkbuf_4 _3939_ (.A(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__o22ai_1 _3940_ (.A1(_0347_),
    .A2(_0349_),
    .B1(_0351_),
    .B2(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__a221oi_1 _3941_ (.A1(_0337_),
    .A2(_0342_),
    .B1(_0343_),
    .B2(_0346_),
    .C1(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__clkbuf_4 _3942_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _3943_ (.A(_3184_),
    .B(_0339_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_2 _3944_ (.A(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__buf_2 _3945_ (.A(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__buf_2 _3946_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _3947_ (.A(_3187_),
    .B(_0339_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_2 _3948_ (.A(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__buf_2 _3949_ (.A(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__inv_2 _3950_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2_2 _3951_ (.A(_3173_),
    .B(_0339_),
    .Y(_0365_));
 sky130_fd_sc_hd__clkbuf_4 _3952_ (.A(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _3953_ (.A(_3178_),
    .B(_0338_),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_2 _3954_ (.A(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__buf_2 _3955_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__buf_2 _3956_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_1 _3957_ (.A(_0369_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__o21ai_1 _3958_ (.A1(_0364_),
    .A2(_0366_),
    .B1(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a221oi_1 _3959_ (.A1(_0356_),
    .A2(_0359_),
    .B1(_0360_),
    .B2(_0363_),
    .C1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _3960_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2_2 _3961_ (.A(_3198_),
    .B(_0339_),
    .Y(_0375_));
 sky130_fd_sc_hd__buf_2 _3962_ (.A(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _3963_ (.A(_3208_),
    .B(_0338_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_2 _3964_ (.A(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__buf_4 _3965_ (.A(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_4 _3966_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_1 _3967_ (.A(_0379_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__and2_1 _3968_ (.A(_3201_),
    .B(_0338_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_2 _3969_ (.A(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_4 _3970_ (.A(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__buf_2 _3971_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _3972_ (.A(_0384_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__inv_2 _3973_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_0387_));
 sky130_fd_sc_hd__nand2_1 _3974_ (.A(_3217_),
    .B(_0339_),
    .Y(_0388_));
 sky130_fd_sc_hd__clkbuf_2 _3975_ (.A(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _3976_ (.A(_0387_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__o2111a_1 _3977_ (.A1(_0374_),
    .A2(_0376_),
    .B1(_0381_),
    .C1(_0386_),
    .D1(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_4 _3978_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _3979_ (.A(_3223_),
    .B(_0338_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_2 _3980_ (.A(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__buf_2 _3981_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__buf_2 _3982_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _3983_ (.A(_3038_),
    .B(_0339_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_2 _3984_ (.A(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_4 _3985_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__and2_1 _3986_ (.A(_3231_),
    .B(_0338_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_2 _3987_ (.A(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__buf_2 _3988_ (.A(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_4 _3989_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_0403_));
 sky130_fd_sc_hd__nand2_1 _3990_ (.A(_0402_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__and2_1 _3991_ (.A(_3237_),
    .B(_0338_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_2 _3992_ (.A(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__buf_2 _3993_ (.A(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_4 _3994_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_0408_));
 sky130_fd_sc_hd__nand2_1 _3995_ (.A(_0407_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_0404_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__a221oi_1 _3997_ (.A1(_0392_),
    .A2(_0395_),
    .B1(_0396_),
    .B2(_0399_),
    .C1(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__and4_1 _3998_ (.A(_0355_),
    .B(_0373_),
    .C(_0391_),
    .D(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__and3_1 _3999_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_4 _4000_ (.A(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _4001_ (.A(_3201_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_2 _4002_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__buf_2 _4003_ (.A(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__and2_1 _4004_ (.A(_3198_),
    .B(_0414_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_2 _4005_ (.A(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__buf_4 _4006_ (.A(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__inv_2 _4007_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_0421_));
 sky130_fd_sc_hd__nand2_2 _4008_ (.A(_3208_),
    .B(_0414_),
    .Y(_0422_));
 sky130_fd_sc_hd__clkbuf_4 _4009_ (.A(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__inv_2 _4010_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_2 _4011_ (.A(_3217_),
    .B(_0414_),
    .Y(_0425_));
 sky130_fd_sc_hd__clkbuf_4 _4012_ (.A(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o22ai_1 _4013_ (.A1(_0421_),
    .A2(_0423_),
    .B1(_0424_),
    .B2(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__a221oi_1 _4014_ (.A1(_3101_),
    .A2(_0417_),
    .B1(_3104_),
    .B2(_0420_),
    .C1(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__and2_1 _4015_ (.A(_3142_),
    .B(_0413_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_2 _4016_ (.A(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__buf_4 _4017_ (.A(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__and2_1 _4018_ (.A(_3151_),
    .B(_0414_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_2 _4019_ (.A(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__buf_6 _4020_ (.A(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__inv_2 _4021_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_0435_));
 sky130_fd_sc_hd__nand2_2 _4022_ (.A(_3164_),
    .B(_0414_),
    .Y(_0436_));
 sky130_fd_sc_hd__buf_2 _4023_ (.A(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__and2_1 _4024_ (.A(_3159_),
    .B(_0413_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_2 _4025_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__buf_2 _4026_ (.A(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__nand2_1 _4027_ (.A(_0440_),
    .B(_3113_),
    .Y(_0441_));
 sky130_fd_sc_hd__o21ai_1 _4028_ (.A1(_0435_),
    .A2(_0437_),
    .B1(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__a221oi_1 _4029_ (.A1(_3107_),
    .A2(_0431_),
    .B1(_3110_),
    .B2(_0434_),
    .C1(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__and2_1 _4030_ (.A(_3184_),
    .B(_0413_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_2 _4031_ (.A(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__buf_2 _4032_ (.A(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__and2_1 _4033_ (.A(_3187_),
    .B(_0414_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_2 _4034_ (.A(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__buf_2 _4035_ (.A(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__inv_2 _4036_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_2 _4037_ (.A(_3173_),
    .B(_0414_),
    .Y(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _4038_ (.A(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__and2_1 _4039_ (.A(_3178_),
    .B(_0413_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_2 _4040_ (.A(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__buf_2 _4041_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__nand2_1 _4042_ (.A(_0455_),
    .B(_3084_),
    .Y(_0456_));
 sky130_fd_sc_hd__o21ai_1 _4043_ (.A1(_0450_),
    .A2(_0452_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__a221oi_1 _4044_ (.A1(_3087_),
    .A2(_0446_),
    .B1(_3090_),
    .B2(_0449_),
    .C1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__and2_1 _4045_ (.A(_3223_),
    .B(_0413_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_2 _4046_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _4047_ (.A(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__and2_1 _4048_ (.A(_3038_),
    .B(_0413_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_2 _4049_ (.A(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_4 _4050_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__inv_2 _4051_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_2 _4052_ (.A(_3237_),
    .B(_0414_),
    .Y(_0466_));
 sky130_fd_sc_hd__buf_2 _4053_ (.A(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__inv_2 _4054_ (.A(_3122_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_2 _4055_ (.A(_3231_),
    .B(_0414_),
    .Y(_0469_));
 sky130_fd_sc_hd__buf_2 _4056_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__o22ai_1 _4057_ (.A1(_0465_),
    .A2(_0467_),
    .B1(_0468_),
    .B2(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__a221oi_1 _4058_ (.A1(_3125_),
    .A2(_0461_),
    .B1(_3129_),
    .B2(_0464_),
    .C1(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__and4_1 _4059_ (.A(_0428_),
    .B(_0443_),
    .C(_0458_),
    .D(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_4 _4060_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_0474_));
 sky130_fd_sc_hd__or3_1 _4061_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .B(_3039_),
    .C(_3248_),
    .X(_0475_));
 sky130_fd_sc_hd__inv_2 _4062_ (.A(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__clkbuf_4 _4063_ (.A(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__and2_1 _4064_ (.A(_3159_),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_2 _4065_ (.A(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__buf_2 _4066_ (.A(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__buf_2 _4067_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_0481_));
 sky130_fd_sc_hd__and2_1 _4068_ (.A(_3164_),
    .B(_0477_),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_2 _4069_ (.A(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__buf_4 _4070_ (.A(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__inv_2 _4071_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_0485_));
 sky130_fd_sc_hd__nand2_2 _4072_ (.A(_3142_),
    .B(_0477_),
    .Y(_0486_));
 sky130_fd_sc_hd__buf_2 _4073_ (.A(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__inv_2 _4074_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_2 _4075_ (.A(_3151_),
    .B(_0477_),
    .Y(_0489_));
 sky130_fd_sc_hd__buf_2 _4076_ (.A(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__o22ai_1 _4077_ (.A1(_0485_),
    .A2(_0487_),
    .B1(_0488_),
    .B2(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__a221oi_1 _4078_ (.A1(_0474_),
    .A2(_0480_),
    .B1(_0481_),
    .B2(_0484_),
    .C1(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _4079_ (.A(_3178_),
    .Y(_0493_));
 sky130_fd_sc_hd__nor2_2 _4080_ (.A(_0475_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__clkbuf_4 _4081_ (.A(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nand2_1 _4082_ (.A(_0495_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_0496_));
 sky130_fd_sc_hd__and2_1 _4083_ (.A(_3187_),
    .B(_0476_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_2 _4084_ (.A(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__buf_2 _4085_ (.A(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__buf_2 _4086_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _4087_ (.A(_0499_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__and2_1 _4088_ (.A(_3173_),
    .B(_0476_),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_2 _4089_ (.A(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__buf_4 _4090_ (.A(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_1 _4091_ (.A(_0504_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_0505_));
 sky130_fd_sc_hd__and2_1 _4092_ (.A(_3184_),
    .B(_0476_),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_2 _4093_ (.A(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__buf_4 _4094_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__nand2_1 _4095_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0509_));
 sky130_fd_sc_hd__and4_1 _4096_ (.A(_0496_),
    .B(_0501_),
    .C(_0505_),
    .D(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__inv_2 _4097_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_2 _4098_ (.A(_3208_),
    .B(_0477_),
    .Y(_0512_));
 sky130_fd_sc_hd__buf_2 _4099_ (.A(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__inv_2 _4100_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_2 _4101_ (.A(_3217_),
    .B(_0477_),
    .Y(_0515_));
 sky130_fd_sc_hd__buf_2 _4102_ (.A(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__o22ai_1 _4103_ (.A1(_0511_),
    .A2(_0513_),
    .B1(_0514_),
    .B2(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__and2_2 _4104_ (.A(_3201_),
    .B(_0477_),
    .X(_0518_));
 sky130_fd_sc_hd__buf_2 _4105_ (.A(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__and2_2 _4106_ (.A(_3198_),
    .B(_0477_),
    .X(_0520_));
 sky130_fd_sc_hd__buf_2 _4107_ (.A(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__buf_2 _4108_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0522_));
 sky130_fd_sc_hd__a22o_1 _4109_ (.A1(_0519_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .B1(_0521_),
    .B2(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__nor2_1 _4110_ (.A(_0517_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__clkbuf_4 _4111_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .X(_0525_));
 sky130_fd_sc_hd__and2_1 _4112_ (.A(_3223_),
    .B(_0476_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_2 _4113_ (.A(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _4114_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__buf_2 _4115_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .X(_0529_));
 sky130_fd_sc_hd__and2_1 _4116_ (.A(_3038_),
    .B(_0476_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_2 _4117_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__buf_2 _4118_ (.A(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__inv_2 _4119_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_2 _4120_ (.A(_3237_),
    .B(_0477_),
    .Y(_0534_));
 sky130_fd_sc_hd__buf_2 _4121_ (.A(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__inv_2 _4122_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_2 _4123_ (.A(_3231_),
    .B(_0477_),
    .Y(_0537_));
 sky130_fd_sc_hd__buf_2 _4124_ (.A(_0537_),
    .X(_0538_));
 sky130_fd_sc_hd__o22ai_1 _4125_ (.A1(_0533_),
    .A2(_0535_),
    .B1(_0536_),
    .B2(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__a221oi_1 _4126_ (.A1(_0525_),
    .A2(_0528_),
    .B1(_0529_),
    .B2(_0532_),
    .C1(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__and4_1 _4127_ (.A(_0492_),
    .B(_0510_),
    .C(_0524_),
    .D(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__buf_2 _4128_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .X(_0542_));
 sky130_fd_sc_hd__or3_1 _4129_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .B(_3039_),
    .C(_3143_),
    .X(_0543_));
 sky130_fd_sc_hd__inv_2 _4130_ (.A(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__buf_2 _4131_ (.A(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _4132_ (.A(_3159_),
    .B(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__clkbuf_2 _4133_ (.A(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__buf_2 _4134_ (.A(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_4 _4135_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .X(_0549_));
 sky130_fd_sc_hd__and2_1 _4136_ (.A(_3164_),
    .B(_0545_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_2 _4137_ (.A(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__buf_4 _4138_ (.A(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__and2_1 _4139_ (.A(_3151_),
    .B(_0545_),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_2 _4140_ (.A(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__buf_6 _4141_ (.A(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _4142_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_1 _4143_ (.A(_0555_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__and2_1 _4144_ (.A(_3142_),
    .B(_0545_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_2 _4145_ (.A(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__buf_4 _4146_ (.A(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__buf_2 _4147_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .X(_0561_));
 sky130_fd_sc_hd__nand2_1 _4148_ (.A(_0560_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(_0557_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__a221oi_1 _4150_ (.A1(_0542_),
    .A2(_0548_),
    .B1(_0549_),
    .B2(_0552_),
    .C1(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__clkbuf_4 _4151_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .X(_0565_));
 sky130_fd_sc_hd__and2_1 _4152_ (.A(_3173_),
    .B(_0545_),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_2 _4153_ (.A(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_4 _4154_ (.A(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__buf_2 _4155_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_2 _4156_ (.A(_0543_),
    .B(_0493_),
    .Y(_0570_));
 sky130_fd_sc_hd__clkbuf_4 _4157_ (.A(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__and2_1 _4158_ (.A(_3187_),
    .B(_0544_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_2 _4159_ (.A(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__buf_2 _4160_ (.A(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__buf_2 _4161_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_1 _4162_ (.A(_0574_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__and2_1 _4163_ (.A(_3184_),
    .B(_0544_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_2 _4164_ (.A(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__buf_4 _4165_ (.A(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__buf_2 _4166_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_1 _4167_ (.A(_0579_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _4168_ (.A(_0576_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__a221oi_1 _4169_ (.A1(_0565_),
    .A2(_0568_),
    .B1(_0569_),
    .B2(_0571_),
    .C1(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__inv_2 _4170_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_0584_));
 sky130_fd_sc_hd__nand2_2 _4171_ (.A(_3198_),
    .B(_0545_),
    .Y(_0585_));
 sky130_fd_sc_hd__buf_2 _4172_ (.A(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__and2_1 _4173_ (.A(_3208_),
    .B(_0544_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_2 _4174_ (.A(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__buf_4 _4175_ (.A(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__buf_2 _4176_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_0590_));
 sky130_fd_sc_hd__nand2_1 _4177_ (.A(_0589_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__and2_1 _4178_ (.A(_3201_),
    .B(_0544_),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_2 _4179_ (.A(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__buf_2 _4180_ (.A(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_4 _4181_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _4182_ (.A(_0594_),
    .B(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _4183_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_2 _4184_ (.A(_3217_),
    .B(_0545_),
    .Y(_0598_));
 sky130_fd_sc_hd__clkbuf_2 _4185_ (.A(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__or2_1 _4186_ (.A(_0597_),
    .B(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__o2111a_1 _4187_ (.A1(_0584_),
    .A2(_0586_),
    .B1(_0591_),
    .C1(_0596_),
    .D1(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__clkbuf_4 _4188_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .X(_0602_));
 sky130_fd_sc_hd__and2_1 _4189_ (.A(_3237_),
    .B(_0545_),
    .X(_0603_));
 sky130_fd_sc_hd__clkbuf_2 _4190_ (.A(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_4 _4191_ (.A(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__clkbuf_4 _4192_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .X(_0606_));
 sky130_fd_sc_hd__and2_1 _4193_ (.A(_3231_),
    .B(_0545_),
    .X(_0607_));
 sky130_fd_sc_hd__clkbuf_2 _4194_ (.A(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_4 _4195_ (.A(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__inv_2 _4196_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_0610_));
 sky130_fd_sc_hd__nand2_2 _4197_ (.A(_3038_),
    .B(_0545_),
    .Y(_0611_));
 sky130_fd_sc_hd__buf_2 _4198_ (.A(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__and2_1 _4199_ (.A(_3223_),
    .B(_0544_),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_2 _4200_ (.A(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__buf_2 _4201_ (.A(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__nand2_1 _4202_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_0616_));
 sky130_fd_sc_hd__o21ai_1 _4203_ (.A1(_0610_),
    .A2(_0612_),
    .B1(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__a221oi_2 _4204_ (.A1(_0602_),
    .A2(_0605_),
    .B1(_0606_),
    .B2(_0609_),
    .C1(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__and4_1 _4205_ (.A(_0564_),
    .B(_0583_),
    .C(_0601_),
    .D(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__and4_1 _4206_ (.A(_0412_),
    .B(_0473_),
    .C(_0541_),
    .D(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__o41a_1 _4207_ (.A1(\egd_top.BitStream_buffer.pc[2] ),
    .A2(\egd_top.BitStream_buffer.pc[3] ),
    .A3(\egd_top.BitStream_buffer.pc[1] ),
    .A4(_3036_),
    .B1(_3250_),
    .X(_0621_));
 sky130_fd_sc_hd__and4b_1 _4208_ (.A_N(_0621_),
    .B(_3039_),
    .C(_3248_),
    .D(_3143_),
    .X(_0622_));
 sky130_fd_sc_hd__clkbuf_2 _4209_ (.A(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__buf_2 _4210_ (.A(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__buf_2 _4211_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0625_));
 sky130_fd_sc_hd__nand2_1 _4212_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand3_1 _4213_ (.A(_0336_),
    .B(_0620_),
    .C(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__nor2_1 _4214_ (.A(_3134_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__nor2_1 _4215_ (.A(_3133_),
    .B(_0628_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21ai_1 _4216_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_0629_));
 sky130_fd_sc_hd__inv_2 _4217_ (.A(_3155_),
    .Y(_0630_));
 sky130_fd_sc_hd__clkbuf_4 _4218_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .X(_0631_));
 sky130_fd_sc_hd__nand2_1 _4219_ (.A(_3154_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__a22o_1 _4220_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_0633_));
 sky130_fd_sc_hd__inv_2 _4221_ (.A(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__o211a_1 _4222_ (.A1(_0630_),
    .A2(_3147_),
    .B1(_0632_),
    .C1(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__inv_2 _4223_ (.A(_3191_),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_1 _4224_ (.A(_3190_),
    .B(_3212_),
    .Y(_0637_));
 sky130_fd_sc_hd__o21ai_1 _4225_ (.A1(_0636_),
    .A2(_3186_),
    .B1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__a221oi_1 _4226_ (.A1(_3177_),
    .A2(_3176_),
    .B1(_3182_),
    .B2(_3181_),
    .C1(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand2_1 _4227_ (.A(_3204_),
    .B(_3195_),
    .Y(_0640_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(_3211_),
    .B(_3214_),
    .Y(_0641_));
 sky130_fd_sc_hd__inv_2 _4229_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .Y(_0642_));
 sky130_fd_sc_hd__or2_1 _4230_ (.A(_0642_),
    .B(_3219_),
    .X(_0643_));
 sky130_fd_sc_hd__o2111a_1 _4231_ (.A1(_3136_),
    .A2(_3200_),
    .B1(_0640_),
    .C1(_0641_),
    .D1(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__nand2_1 _4232_ (.A(_3234_),
    .B(_3222_),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _4233_ (.A(_3240_),
    .B(_3235_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _4234_ (.A(_0645_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__a221oi_1 _4235_ (.A1(_3227_),
    .A2(_3226_),
    .B1(_3351_),
    .B2(_3230_),
    .C1(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__and4_1 _4236_ (.A(_0635_),
    .B(_0639_),
    .C(_0644_),
    .D(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__inv_2 _4237_ (.A(_3256_),
    .Y(_0650_));
 sky130_fd_sc_hd__nand2_1 _4238_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_0651_));
 sky130_fd_sc_hd__nand2_1 _4239_ (.A(_3260_),
    .B(_3246_),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _4240_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0653_));
 sky130_fd_sc_hd__or2_1 _4241_ (.A(_0653_),
    .B(_3265_),
    .X(_0654_));
 sky130_fd_sc_hd__o2111a_1 _4242_ (.A1(_0650_),
    .A2(_3252_),
    .B1(_0651_),
    .C1(_0652_),
    .D1(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(_3273_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _4244_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_0657_));
 sky130_fd_sc_hd__inv_2 _4245_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0658_));
 sky130_fd_sc_hd__or2_1 _4246_ (.A(_0658_),
    .B(_3281_),
    .X(_0659_));
 sky130_fd_sc_hd__o2111a_1 _4247_ (.A1(_3303_),
    .A2(_3270_),
    .B1(_0656_),
    .C1(_0657_),
    .D1(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__inv_2 _4248_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0661_));
 sky130_fd_sc_hd__or2_1 _4249_ (.A(_0661_),
    .B(_3294_),
    .X(_0662_));
 sky130_fd_sc_hd__o221a_1 _4250_ (.A1(_3292_),
    .A2(_3287_),
    .B1(_3285_),
    .B2(_3290_),
    .C1(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__inv_2 _4251_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_0664_));
 sky130_fd_sc_hd__o22ai_1 _4252_ (.A1(_3306_),
    .A2(_3305_),
    .B1(_0664_),
    .B2(_3308_),
    .Y(_0665_));
 sky130_fd_sc_hd__a221oi_1 _4253_ (.A1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .A2(_3299_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .B2(_3302_),
    .C1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__and4_1 _4254_ (.A(_0655_),
    .B(_0660_),
    .C(_0663_),
    .D(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__inv_2 _4255_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .Y(_0668_));
 sky130_fd_sc_hd__o22ai_1 _4256_ (.A1(_3326_),
    .A2(_3324_),
    .B1(_0668_),
    .B2(_3328_),
    .Y(_0669_));
 sky130_fd_sc_hd__a221oi_1 _4257_ (.A1(_3318_),
    .A2(_3317_),
    .B1(_3347_),
    .B2(_3321_),
    .C1(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _4258_ (.A(_3341_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _4259_ (.A(_3346_),
    .B(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2_1 _4260_ (.A(_0671_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__a221oi_1 _4261_ (.A1(_3335_),
    .A2(_3334_),
    .B1(_3369_),
    .B2(_3338_),
    .C1(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__buf_2 _4262_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_0675_));
 sky130_fd_sc_hd__inv_2 _4263_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_0676_));
 sky130_fd_sc_hd__buf_2 _4264_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_0677_));
 sky130_fd_sc_hd__nand2_1 _4265_ (.A(_3364_),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__o21ai_1 _4266_ (.A1(_0676_),
    .A2(_3361_),
    .B1(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__a221oi_1 _4267_ (.A1(_3355_),
    .A2(_3354_),
    .B1(_0675_),
    .B2(_3358_),
    .C1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__buf_2 _4268_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_1 _4269_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_0682_));
 sky130_fd_sc_hd__o21ai_1 _4270_ (.A1(_3431_),
    .A2(_3379_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__a221oi_1 _4271_ (.A1(_3373_),
    .A2(_3372_),
    .B1(_0681_),
    .B2(_3376_),
    .C1(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__and4_1 _4272_ (.A(_0670_),
    .B(_0674_),
    .C(_0680_),
    .D(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__inv_2 _4273_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0686_));
 sky130_fd_sc_hd__buf_2 _4274_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .X(_0687_));
 sky130_fd_sc_hd__nand2_1 _4275_ (.A(_3393_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__buf_2 _4276_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_1 _4277_ (.A(_3398_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__inv_2 _4278_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0691_));
 sky130_fd_sc_hd__or2_1 _4279_ (.A(_0691_),
    .B(_3403_),
    .X(_0692_));
 sky130_fd_sc_hd__o2111a_1 _4280_ (.A1(_0686_),
    .A2(_3390_),
    .B1(_0688_),
    .C1(_0690_),
    .D1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__inv_2 _4281_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .Y(_0694_));
 sky130_fd_sc_hd__nand2_1 _4282_ (.A(_3411_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0695_));
 sky130_fd_sc_hd__buf_2 _4283_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_3415_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__inv_2 _4285_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0698_));
 sky130_fd_sc_hd__or2_1 _4286_ (.A(_0698_),
    .B(_3420_),
    .X(_0699_));
 sky130_fd_sc_hd__o2111a_1 _4287_ (.A1(_0694_),
    .A2(_3408_),
    .B1(_0695_),
    .C1(_0697_),
    .D1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__inv_2 _4288_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _4289_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_0702_));
 sky130_fd_sc_hd__o21ai_1 _4290_ (.A1(_0701_),
    .A2(_3433_),
    .B1(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__a221oi_1 _4291_ (.A1(_3427_),
    .A2(_3426_),
    .B1(_3399_),
    .B2(_3430_),
    .C1(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__buf_2 _4292_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .X(_0705_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(_0331_),
    .B(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_0706_));
 sky130_fd_sc_hd__o21ai_1 _4294_ (.A1(_0364_),
    .A2(_0328_),
    .B1(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__a221oi_1 _4295_ (.A1(_0322_),
    .A2(_3443_),
    .B1(_0705_),
    .B2(_0325_),
    .C1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__and4_1 _4296_ (.A(_0693_),
    .B(_0700_),
    .C(_0704_),
    .D(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__and4_1 _4297_ (.A(_0649_),
    .B(_0667_),
    .C(_0685_),
    .D(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__inv_2 _4298_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_0711_));
 sky130_fd_sc_hd__o22ai_1 _4299_ (.A1(_0351_),
    .A2(_0349_),
    .B1(_0711_),
    .B2(_0353_),
    .Y(_0712_));
 sky130_fd_sc_hd__a221oi_1 _4300_ (.A1(_0343_),
    .A2(_0342_),
    .B1(_0408_),
    .B2(_0346_),
    .C1(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__inv_2 _4301_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_0714_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_0369_),
    .B(_0356_),
    .Y(_0715_));
 sky130_fd_sc_hd__o21ai_1 _4303_ (.A1(_0714_),
    .A2(_0366_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a221oi_1 _4304_ (.A1(_0360_),
    .A2(_0359_),
    .B1(_0380_),
    .B2(_0363_),
    .C1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__buf_2 _4305_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_0718_));
 sky130_fd_sc_hd__nand2_1 _4306_ (.A(_0379_),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__buf_2 _4307_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_0720_));
 sky130_fd_sc_hd__nand2_1 _4308_ (.A(_0384_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__inv_2 _4309_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_0722_));
 sky130_fd_sc_hd__or2_1 _4310_ (.A(_0722_),
    .B(_0389_),
    .X(_0723_));
 sky130_fd_sc_hd__o2111a_1 _4311_ (.A1(_0347_),
    .A2(_0376_),
    .B1(_0719_),
    .C1(_0721_),
    .D1(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__buf_2 _4312_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_0725_));
 sky130_fd_sc_hd__nand2_1 _4313_ (.A(_0402_),
    .B(_0392_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_0407_),
    .B(_0403_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _4315_ (.A(_0726_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__a221oi_1 _4316_ (.A1(_0396_),
    .A2(_0395_),
    .B1(_0725_),
    .B2(_0399_),
    .C1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__and4_1 _4317_ (.A(_0713_),
    .B(_0717_),
    .C(_0724_),
    .D(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__inv_2 _4318_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_0731_));
 sky130_fd_sc_hd__o22ai_1 _4319_ (.A1(_0424_),
    .A2(_0423_),
    .B1(_0731_),
    .B2(_0426_),
    .Y(_0732_));
 sky130_fd_sc_hd__a221oi_1 _4320_ (.A1(_3104_),
    .A2(_0417_),
    .B1(_3107_),
    .B2(_0420_),
    .C1(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _4321_ (.A(_0440_),
    .B(_3116_),
    .Y(_0734_));
 sky130_fd_sc_hd__o21ai_1 _4322_ (.A1(_0465_),
    .A2(_0437_),
    .B1(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__a221oi_1 _4323_ (.A1(_3110_),
    .A2(_0431_),
    .B1(_3113_),
    .B2(_0434_),
    .C1(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__inv_2 _4324_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(_0455_),
    .B(_3087_),
    .Y(_0738_));
 sky130_fd_sc_hd__o21ai_1 _4326_ (.A1(_0737_),
    .A2(_0452_),
    .B1(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__a221oi_1 _4327_ (.A1(_3090_),
    .A2(_0446_),
    .B1(_3093_),
    .B2(_0449_),
    .C1(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__inv_2 _4328_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_0741_));
 sky130_fd_sc_hd__o22ai_1 _4329_ (.A1(_0468_),
    .A2(_0467_),
    .B1(_0741_),
    .B2(_0470_),
    .Y(_0742_));
 sky130_fd_sc_hd__a221oi_1 _4330_ (.A1(_3129_),
    .A2(_0461_),
    .B1(_0625_),
    .B2(_0464_),
    .C1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__and4_1 _4331_ (.A(_0733_),
    .B(_0736_),
    .C(_0740_),
    .D(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__buf_2 _4332_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_0745_));
 sky130_fd_sc_hd__inv_2 _4333_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_0746_));
 sky130_fd_sc_hd__o22ai_1 _4334_ (.A1(_0488_),
    .A2(_0487_),
    .B1(_0746_),
    .B2(_0490_),
    .Y(_0747_));
 sky130_fd_sc_hd__a221oi_1 _4335_ (.A1(_0481_),
    .A2(_0480_),
    .B1(_0745_),
    .B2(_0484_),
    .C1(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__buf_2 _4336_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .X(_0749_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_0495_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__buf_2 _4338_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .X(_0751_));
 sky130_fd_sc_hd__nand2_1 _4339_ (.A(_0499_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _4340_ (.A(_0504_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_1 _4341_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0754_));
 sky130_fd_sc_hd__and4_1 _4342_ (.A(_0750_),
    .B(_0752_),
    .C(_0753_),
    .D(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__inv_2 _4343_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0756_));
 sky130_fd_sc_hd__o22ai_1 _4344_ (.A1(_0514_),
    .A2(_0513_),
    .B1(_0756_),
    .B2(_0516_),
    .Y(_0757_));
 sky130_fd_sc_hd__clkbuf_4 _4345_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_0758_));
 sky130_fd_sc_hd__a22o_1 _4346_ (.A1(_0519_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .B1(_0521_),
    .B2(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nor2_1 _4347_ (.A(_0757_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__inv_2 _4348_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_0761_));
 sky130_fd_sc_hd__o22ai_1 _4349_ (.A1(_0536_),
    .A2(_0535_),
    .B1(_0761_),
    .B2(_0538_),
    .Y(_0762_));
 sky130_fd_sc_hd__a221oi_1 _4350_ (.A1(_0529_),
    .A2(_0528_),
    .B1(_0565_),
    .B2(_0532_),
    .C1(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__and4_1 _4351_ (.A(_0748_),
    .B(_0755_),
    .C(_0760_),
    .D(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__nand2_1 _4352_ (.A(_0555_),
    .B(_0542_),
    .Y(_0765_));
 sky130_fd_sc_hd__nand2_1 _4353_ (.A(_0560_),
    .B(_0556_),
    .Y(_0766_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_0765_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__a221oi_1 _4355_ (.A1(_0549_),
    .A2(_0548_),
    .B1(_0602_),
    .B2(_0552_),
    .C1(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__nand2_1 _4356_ (.A(_0574_),
    .B(_0590_),
    .Y(_0769_));
 sky130_fd_sc_hd__nand2_1 _4357_ (.A(_0579_),
    .B(_0575_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _4358_ (.A(_0769_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__a221oi_1 _4359_ (.A1(_0569_),
    .A2(_0568_),
    .B1(_0580_),
    .B2(_0571_),
    .C1(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__inv_2 _4360_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0773_));
 sky130_fd_sc_hd__clkbuf_4 _4361_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _4362_ (.A(_0589_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__buf_2 _4363_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_0776_));
 sky130_fd_sc_hd__nand2_1 _4364_ (.A(_0594_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_2 _4365_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_0778_));
 sky130_fd_sc_hd__or2_1 _4366_ (.A(_0778_),
    .B(_0599_),
    .X(_0779_));
 sky130_fd_sc_hd__o2111a_1 _4367_ (.A1(_0773_),
    .A2(_0586_),
    .B1(_0775_),
    .C1(_0777_),
    .D1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__buf_2 _4368_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _4369_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_0782_));
 sky130_fd_sc_hd__o21ai_1 _4370_ (.A1(_0450_),
    .A2(_0612_),
    .B1(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__a221oi_1 _4371_ (.A1(_0606_),
    .A2(_0605_),
    .B1(_0781_),
    .B2(_0609_),
    .C1(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__and4_1 _4372_ (.A(_0768_),
    .B(_0772_),
    .C(_0780_),
    .D(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__and4_1 _4373_ (.A(_0730_),
    .B(_0744_),
    .C(_0764_),
    .D(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__buf_2 _4374_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0787_));
 sky130_fd_sc_hd__nand2_1 _4375_ (.A(_0624_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__nand3_1 _4376_ (.A(_0710_),
    .B(_0786_),
    .C(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__nor2_1 _4377_ (.A(_3134_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_1 _4378_ (.A(_0629_),
    .B(_0790_),
    .Y(_0296_));
 sky130_fd_sc_hd__o21ai_1 _4379_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_0791_));
 sky130_fd_sc_hd__inv_2 _4380_ (.A(_0631_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_1 _4381_ (.A(_3154_),
    .B(_3167_),
    .Y(_0793_));
 sky130_fd_sc_hd__a22o_1 _4382_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_0794_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__o211a_1 _4384_ (.A1(_0792_),
    .A2(_3147_),
    .B1(_0793_),
    .C1(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__inv_2 _4385_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .Y(_0797_));
 sky130_fd_sc_hd__nand2_1 _4386_ (.A(_3190_),
    .B(_3214_),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_1 _4387_ (.A1(_0797_),
    .A2(_3186_),
    .B1(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__a221oi_1 _4388_ (.A1(_3182_),
    .A2(_3176_),
    .B1(_3191_),
    .B2(_3181_),
    .C1(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_3204_),
    .B(_3135_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_1 _4390_ (.A(_3211_),
    .B(_3205_),
    .Y(_0802_));
 sky130_fd_sc_hd__or2_1 _4391_ (.A(_3196_),
    .B(_3219_),
    .X(_0803_));
 sky130_fd_sc_hd__o2111a_1 _4392_ (.A1(_0630_),
    .A2(_3200_),
    .B1(_0801_),
    .C1(_0802_),
    .D1(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__nand2_1 _4393_ (.A(_3234_),
    .B(_3227_),
    .Y(_0805_));
 sky130_fd_sc_hd__nand2_1 _4394_ (.A(_3240_),
    .B(_3222_),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2_1 _4395_ (.A(_0805_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__a221oi_1 _4396_ (.A1(_3351_),
    .A2(_3226_),
    .B1(_3355_),
    .B2(_3230_),
    .C1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__and4_1 _4397_ (.A(_0796_),
    .B(_0800_),
    .C(_0804_),
    .D(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__nand2_1 _4398_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _4399_ (.A(_3260_),
    .B(_3256_),
    .Y(_0811_));
 sky130_fd_sc_hd__or2_1 _4400_ (.A(_3279_),
    .B(_3265_),
    .X(_0812_));
 sky130_fd_sc_hd__o2111a_1 _4401_ (.A1(_3263_),
    .A2(_3252_),
    .B1(_0810_),
    .C1(_0811_),
    .D1(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__nand2_1 _4402_ (.A(_3273_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0814_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0815_));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(_3268_),
    .B(_3281_),
    .X(_0816_));
 sky130_fd_sc_hd__o2111a_1 _4405_ (.A1(_3306_),
    .A2(_3270_),
    .B1(_0814_),
    .C1(_0815_),
    .D1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__or2_1 _4406_ (.A(_3247_),
    .B(_3294_),
    .X(_0818_));
 sky130_fd_sc_hd__o221a_1 _4407_ (.A1(_0661_),
    .A2(_3287_),
    .B1(_3292_),
    .B2(_3290_),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__inv_2 _4408_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_0820_));
 sky130_fd_sc_hd__o22ai_1 _4409_ (.A1(_0664_),
    .A2(_3305_),
    .B1(_0820_),
    .B2(_3308_),
    .Y(_0821_));
 sky130_fd_sc_hd__a221oi_1 _4410_ (.A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .A2(_3299_),
    .B1(_3177_),
    .B2(_3302_),
    .C1(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__and4_1 _4411_ (.A(_0813_),
    .B(_0817_),
    .C(_0819_),
    .D(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__inv_2 _4412_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_0824_));
 sky130_fd_sc_hd__o22ai_1 _4413_ (.A1(_0668_),
    .A2(_3324_),
    .B1(_0824_),
    .B2(_3328_),
    .Y(_0825_));
 sky130_fd_sc_hd__a221oi_1 _4414_ (.A1(_3347_),
    .A2(_3317_),
    .B1(_3342_),
    .B2(_3321_),
    .C1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand2_1 _4415_ (.A(_3341_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_0827_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(_3346_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _4417_ (.A(_0827_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__a221oi_1 _4418_ (.A1(_3369_),
    .A2(_3334_),
    .B1(_3373_),
    .B2(_3338_),
    .C1(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_3364_),
    .B(_3325_),
    .Y(_0831_));
 sky130_fd_sc_hd__o21ai_1 _4420_ (.A1(_3322_),
    .A2(_3361_),
    .B1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__a221oi_1 _4421_ (.A1(_0675_),
    .A2(_3354_),
    .B1(_3365_),
    .B2(_3358_),
    .C1(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__buf_2 _4422_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_0834_));
 sky130_fd_sc_hd__nand2_1 _4423_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .Y(_0835_));
 sky130_fd_sc_hd__o21ai_1 _4424_ (.A1(_0701_),
    .A2(_3379_),
    .B1(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__a221oi_1 _4425_ (.A1(_0681_),
    .A2(_3372_),
    .B1(_0834_),
    .B2(_3376_),
    .C1(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__and4_1 _4426_ (.A(_0826_),
    .B(_0830_),
    .C(_0833_),
    .D(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_2 _4427_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .X(_0839_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(_3393_),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__nand2_1 _4429_ (.A(_3398_),
    .B(_3394_),
    .Y(_0841_));
 sky130_fd_sc_hd__or2_1 _4430_ (.A(_3418_),
    .B(_3403_),
    .X(_0842_));
 sky130_fd_sc_hd__o2111a_1 _4431_ (.A1(_3401_),
    .A2(_3390_),
    .B1(_0840_),
    .C1(_0841_),
    .D1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__inv_2 _4432_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .Y(_0844_));
 sky130_fd_sc_hd__nand2_1 _4433_ (.A(_3411_),
    .B(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _4434_ (.A(_3415_),
    .B(_3440_),
    .Y(_0846_));
 sky130_fd_sc_hd__or2_1 _4435_ (.A(_3406_),
    .B(_3420_),
    .X(_0847_));
 sky130_fd_sc_hd__o2111a_1 _4436_ (.A1(_0844_),
    .A2(_3408_),
    .B1(_0845_),
    .C1(_0846_),
    .D1(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__inv_2 _4437_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_0850_));
 sky130_fd_sc_hd__o21ai_1 _4439_ (.A1(_0849_),
    .A2(_3433_),
    .B1(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__a221oi_1 _4440_ (.A1(_3399_),
    .A2(_3426_),
    .B1(_0689_),
    .B2(_3430_),
    .C1(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__buf_2 _4441_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .X(_0853_));
 sky130_fd_sc_hd__buf_2 _4442_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _4443_ (.A(_0331_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__o21ai_1 _4444_ (.A1(_0714_),
    .A2(_0328_),
    .B1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__a221oi_1 _4445_ (.A1(_0705_),
    .A2(_3443_),
    .B1(_0853_),
    .B2(_0325_),
    .C1(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__and4_1 _4446_ (.A(_0843_),
    .B(_0848_),
    .C(_0852_),
    .D(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__and4_1 _4447_ (.A(_0809_),
    .B(_0823_),
    .C(_0838_),
    .D(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__inv_2 _4448_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_0860_));
 sky130_fd_sc_hd__o22ai_1 _4449_ (.A1(_0711_),
    .A2(_0349_),
    .B1(_0860_),
    .B2(_0353_),
    .Y(_0861_));
 sky130_fd_sc_hd__a221oi_1 _4450_ (.A1(_0408_),
    .A2(_0342_),
    .B1(_0403_),
    .B2(_0346_),
    .C1(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__inv_2 _4451_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_0863_));
 sky130_fd_sc_hd__nand2_1 _4452_ (.A(_0369_),
    .B(_0360_),
    .Y(_0864_));
 sky130_fd_sc_hd__o21ai_1 _4453_ (.A1(_0863_),
    .A2(_0366_),
    .B1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__a221oi_1 _4454_ (.A1(_0380_),
    .A2(_0359_),
    .B1(_0718_),
    .B2(_0363_),
    .C1(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand2_1 _4455_ (.A(_0379_),
    .B(_0385_),
    .Y(_0867_));
 sky130_fd_sc_hd__buf_2 _4456_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_0868_));
 sky130_fd_sc_hd__nand2_1 _4457_ (.A(_0384_),
    .B(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__or2_1 _4458_ (.A(_0374_),
    .B(_0389_),
    .X(_0870_));
 sky130_fd_sc_hd__o2111a_1 _4459_ (.A1(_0351_),
    .A2(_0376_),
    .B1(_0867_),
    .C1(_0869_),
    .D1(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__clkbuf_4 _4460_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .X(_0872_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_0402_),
    .B(_0396_),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(_0407_),
    .B(_0392_),
    .Y(_0874_));
 sky130_fd_sc_hd__nand2_1 _4463_ (.A(_0873_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__a221oi_1 _4464_ (.A1(_0725_),
    .A2(_0395_),
    .B1(_0872_),
    .B2(_0399_),
    .C1(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__and4_1 _4465_ (.A(_0862_),
    .B(_0866_),
    .C(_0871_),
    .D(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__inv_2 _4466_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_0878_));
 sky130_fd_sc_hd__o22ai_1 _4467_ (.A1(_0731_),
    .A2(_0423_),
    .B1(_0878_),
    .B2(_0426_),
    .Y(_0879_));
 sky130_fd_sc_hd__a221oi_1 _4468_ (.A1(_3107_),
    .A2(_0417_),
    .B1(_3110_),
    .B2(_0420_),
    .C1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _4469_ (.A(_0440_),
    .B(_3119_),
    .Y(_0881_));
 sky130_fd_sc_hd__o21ai_1 _4470_ (.A1(_0468_),
    .A2(_0437_),
    .B1(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__a221oi_1 _4471_ (.A1(_3113_),
    .A2(_0431_),
    .B1(_3116_),
    .B2(_0434_),
    .C1(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__inv_2 _4472_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_0884_));
 sky130_fd_sc_hd__nand2_1 _4473_ (.A(_0455_),
    .B(_3090_),
    .Y(_0885_));
 sky130_fd_sc_hd__o21ai_1 _4474_ (.A1(_0884_),
    .A2(_0452_),
    .B1(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__a221oi_1 _4475_ (.A1(_3093_),
    .A2(_0446_),
    .B1(_3098_),
    .B2(_0449_),
    .C1(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_2 _4476_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_0888_));
 sky130_fd_sc_hd__o22ai_1 _4477_ (.A1(_0741_),
    .A2(_0467_),
    .B1(_0888_),
    .B2(_0470_),
    .Y(_0889_));
 sky130_fd_sc_hd__a221oi_1 _4478_ (.A1(_0625_),
    .A2(_0461_),
    .B1(_0787_),
    .B2(_0464_),
    .C1(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__and4_1 _4479_ (.A(_0880_),
    .B(_0883_),
    .C(_0887_),
    .D(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_4 _4480_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0892_));
 sky130_fd_sc_hd__inv_2 _4481_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_0893_));
 sky130_fd_sc_hd__o22ai_1 _4482_ (.A1(_0746_),
    .A2(_0487_),
    .B1(_0893_),
    .B2(_0490_),
    .Y(_0894_));
 sky130_fd_sc_hd__a221oi_1 _4483_ (.A1(_0745_),
    .A2(_0480_),
    .B1(_0892_),
    .B2(_0484_),
    .C1(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand2_1 _4484_ (.A(_0495_),
    .B(_0500_),
    .Y(_0896_));
 sky130_fd_sc_hd__buf_2 _4485_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _4486_ (.A(_0499_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_1 _4487_ (.A(_0504_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _4488_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0900_));
 sky130_fd_sc_hd__and4_1 _4489_ (.A(_0896_),
    .B(_0898_),
    .C(_0899_),
    .D(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__inv_2 _4490_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_0902_));
 sky130_fd_sc_hd__o22ai_1 _4491_ (.A1(_0756_),
    .A2(_0513_),
    .B1(_0902_),
    .B2(_0516_),
    .Y(_0903_));
 sky130_fd_sc_hd__clkbuf_4 _4492_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _4493_ (.A1(_0519_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .B1(_0521_),
    .B2(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_1 _4494_ (.A(_0903_),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__inv_2 _4495_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_0907_));
 sky130_fd_sc_hd__o22ai_1 _4496_ (.A1(_0761_),
    .A2(_0535_),
    .B1(_0907_),
    .B2(_0538_),
    .Y(_0908_));
 sky130_fd_sc_hd__a221oi_1 _4497_ (.A1(_0565_),
    .A2(_0528_),
    .B1(_0569_),
    .B2(_0532_),
    .C1(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__and4_1 _4498_ (.A(_0895_),
    .B(_0901_),
    .C(_0906_),
    .D(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_0555_),
    .B(_0549_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _4500_ (.A(_0560_),
    .B(_0542_),
    .Y(_0912_));
 sky130_fd_sc_hd__nand2_1 _4501_ (.A(_0911_),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__a221oi_1 _4502_ (.A1(_0602_),
    .A2(_0548_),
    .B1(_0606_),
    .B2(_0552_),
    .C1(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand2_1 _4503_ (.A(_0574_),
    .B(_0774_),
    .Y(_0915_));
 sky130_fd_sc_hd__nand2_1 _4504_ (.A(_0579_),
    .B(_0590_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_1 _4505_ (.A(_0915_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a221oi_1 _4506_ (.A1(_0580_),
    .A2(_0568_),
    .B1(_0575_),
    .B2(_0571_),
    .C1(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__inv_2 _4507_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_0919_));
 sky130_fd_sc_hd__nand2_1 _4508_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_0920_));
 sky130_fd_sc_hd__nand2_1 _4509_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0921_));
 sky130_fd_sc_hd__or2_1 _4510_ (.A(_0584_),
    .B(_0599_),
    .X(_0922_));
 sky130_fd_sc_hd__o2111a_1 _4511_ (.A1(_0919_),
    .A2(_0586_),
    .B1(_0920_),
    .C1(_0921_),
    .D1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_4 _4512_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .X(_0924_));
 sky130_fd_sc_hd__nand2_1 _4513_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_0925_));
 sky130_fd_sc_hd__o21ai_1 _4514_ (.A1(_0737_),
    .A2(_0612_),
    .B1(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__a221oi_1 _4515_ (.A1(_0781_),
    .A2(_0605_),
    .B1(_0924_),
    .B2(_0609_),
    .C1(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__and4_1 _4516_ (.A(_0914_),
    .B(_0918_),
    .C(_0923_),
    .D(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__and4_1 _4517_ (.A(_0877_),
    .B(_0891_),
    .C(_0910_),
    .D(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__nand2_1 _4518_ (.A(_0624_),
    .B(_3284_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand3_1 _4519_ (.A(_0859_),
    .B(_0929_),
    .C(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__nor2_1 _4520_ (.A(_3134_),
    .B(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__nor2_1 _4521_ (.A(_0791_),
    .B(_0932_),
    .Y(_0295_));
 sky130_fd_sc_hd__o21ai_1 _4522_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_0933_));
 sky130_fd_sc_hd__inv_2 _4523_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_3154_),
    .B(_3241_),
    .Y(_0935_));
 sky130_fd_sc_hd__a22o_1 _4525_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_0936_));
 sky130_fd_sc_hd__inv_2 _4526_ (.A(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__o211a_1 _4527_ (.A1(_0934_),
    .A2(_3147_),
    .B1(_0935_),
    .C1(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__nand2_1 _4528_ (.A(_3190_),
    .B(_3205_),
    .Y(_0939_));
 sky130_fd_sc_hd__o21ai_1 _4529_ (.A1(_3215_),
    .A2(_3186_),
    .B1(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__a221oi_1 _4530_ (.A1(_3191_),
    .A2(_3176_),
    .B1(_3212_),
    .B2(_3181_),
    .C1(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__nand2_1 _4531_ (.A(_3204_),
    .B(_3155_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _4532_ (.A(_3211_),
    .B(_3195_),
    .Y(_0943_));
 sky130_fd_sc_hd__or2_1 _4533_ (.A(_3136_),
    .B(_3219_),
    .X(_0944_));
 sky130_fd_sc_hd__o2111a_1 _4534_ (.A1(_0792_),
    .A2(_3200_),
    .B1(_0942_),
    .C1(_0943_),
    .D1(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__nand2_1 _4535_ (.A(_3234_),
    .B(_3351_),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(_3240_),
    .B(_3227_),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _4537_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__a221oi_1 _4538_ (.A1(_3355_),
    .A2(_3226_),
    .B1(_0675_),
    .B2(_3230_),
    .C1(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__and4_1 _4539_ (.A(_0938_),
    .B(_0941_),
    .C(_0945_),
    .D(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__nand2_1 _4540_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _4541_ (.A(_3260_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_0952_));
 sky130_fd_sc_hd__or2_1 _4542_ (.A(_0658_),
    .B(_3265_),
    .X(_0953_));
 sky130_fd_sc_hd__o2111a_1 _4543_ (.A1(_0653_),
    .A2(_3252_),
    .B1(_0951_),
    .C1(_0952_),
    .D1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__nand2_1 _4544_ (.A(_3273_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _4545_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_0956_));
 sky130_fd_sc_hd__or2_1 _4546_ (.A(_3303_),
    .B(_3281_),
    .X(_0957_));
 sky130_fd_sc_hd__o2111a_1 _4547_ (.A1(_0664_),
    .A2(_3270_),
    .B1(_0955_),
    .C1(_0956_),
    .D1(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__or2_1 _4548_ (.A(_0650_),
    .B(_3294_),
    .X(_0959_));
 sky130_fd_sc_hd__o221a_1 _4549_ (.A1(_3247_),
    .A2(_3287_),
    .B1(_0661_),
    .B2(_3290_),
    .C1(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__inv_2 _4550_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_0961_));
 sky130_fd_sc_hd__o22ai_1 _4551_ (.A1(_0820_),
    .A2(_3305_),
    .B1(_0961_),
    .B2(_3308_),
    .Y(_0962_));
 sky130_fd_sc_hd__a221oi_1 _4552_ (.A1(_3177_),
    .A2(_3299_),
    .B1(_3182_),
    .B2(_3302_),
    .C1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__and4_1 _4553_ (.A(_0954_),
    .B(_0958_),
    .C(_0960_),
    .D(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__inv_2 _4554_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_0965_));
 sky130_fd_sc_hd__o22ai_1 _4555_ (.A1(_0824_),
    .A2(_3324_),
    .B1(_0965_),
    .B2(_3328_),
    .Y(_0966_));
 sky130_fd_sc_hd__a221oi_1 _4556_ (.A1(_3342_),
    .A2(_3317_),
    .B1(_3331_),
    .B2(_3321_),
    .C1(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_3341_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_0968_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_3346_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_0969_));
 sky130_fd_sc_hd__nand2_1 _4559_ (.A(_0968_),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__a221oi_1 _4560_ (.A1(_3373_),
    .A2(_3334_),
    .B1(_0681_),
    .B2(_3338_),
    .C1(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_3364_),
    .B(_3312_),
    .Y(_0972_));
 sky130_fd_sc_hd__o21ai_1 _4562_ (.A1(_3326_),
    .A2(_3361_),
    .B1(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__a221oi_1 _4563_ (.A1(_3365_),
    .A2(_3354_),
    .B1(_0677_),
    .B2(_3358_),
    .C1(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__buf_2 _4564_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .X(_0975_));
 sky130_fd_sc_hd__nand2_1 _4565_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_0976_));
 sky130_fd_sc_hd__o21ai_1 _4566_ (.A1(_0849_),
    .A2(_3379_),
    .B1(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__a221oi_1 _4567_ (.A1(_0834_),
    .A2(_3372_),
    .B1(_0975_),
    .B2(_3376_),
    .C1(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__and4_1 _4568_ (.A(_0967_),
    .B(_0971_),
    .C(_0974_),
    .D(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__buf_2 _4569_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .X(_0980_));
 sky130_fd_sc_hd__nand2_1 _4570_ (.A(_3393_),
    .B(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__nand2_1 _4571_ (.A(_3398_),
    .B(_0687_),
    .Y(_0982_));
 sky130_fd_sc_hd__or2_1 _4572_ (.A(_0698_),
    .B(_3403_),
    .X(_0983_));
 sky130_fd_sc_hd__o2111a_1 _4573_ (.A1(_0691_),
    .A2(_3390_),
    .B1(_0981_),
    .C1(_0982_),
    .D1(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__inv_2 _4574_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_0985_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_3411_),
    .B(_0696_),
    .Y(_0986_));
 sky130_fd_sc_hd__nand2_1 _4576_ (.A(_3415_),
    .B(_0322_),
    .Y(_0987_));
 sky130_fd_sc_hd__or2_1 _4577_ (.A(_0694_),
    .B(_3420_),
    .X(_0988_));
 sky130_fd_sc_hd__o2111a_1 _4578_ (.A1(_0985_),
    .A2(_3408_),
    .B1(_0986_),
    .C1(_0987_),
    .D1(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__inv_2 _4579_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_0990_));
 sky130_fd_sc_hd__nand2_1 _4580_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_0991_));
 sky130_fd_sc_hd__o21ai_1 _4581_ (.A1(_0990_),
    .A2(_3433_),
    .B1(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__a221oi_1 _4582_ (.A1(_0689_),
    .A2(_3426_),
    .B1(_3394_),
    .B2(_3430_),
    .C1(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__nand2_1 _4583_ (.A(_0331_),
    .B(_0370_),
    .Y(_0994_));
 sky130_fd_sc_hd__o21ai_1 _4584_ (.A1(_0863_),
    .A2(_0328_),
    .B1(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__a221oi_1 _4585_ (.A1(_0853_),
    .A2(_3443_),
    .B1(_0854_),
    .B2(_0325_),
    .C1(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__and4_1 _4586_ (.A(_0984_),
    .B(_0989_),
    .C(_0993_),
    .D(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__and4_1 _4587_ (.A(_0950_),
    .B(_0964_),
    .C(_0979_),
    .D(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__inv_2 _4588_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_0999_));
 sky130_fd_sc_hd__o22ai_1 _4589_ (.A1(_0860_),
    .A2(_0349_),
    .B1(_0999_),
    .B2(_0353_),
    .Y(_1000_));
 sky130_fd_sc_hd__a221oi_1 _4590_ (.A1(_0403_),
    .A2(_0342_),
    .B1(_0392_),
    .B2(_0346_),
    .C1(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__inv_2 _4591_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_1002_));
 sky130_fd_sc_hd__nand2_1 _4592_ (.A(_0369_),
    .B(_0380_),
    .Y(_1003_));
 sky130_fd_sc_hd__o21ai_1 _4593_ (.A1(_1002_),
    .A2(_0366_),
    .B1(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__a221oi_1 _4594_ (.A1(_0718_),
    .A2(_0359_),
    .B1(_0385_),
    .B2(_0363_),
    .C1(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__nand2_1 _4595_ (.A(_0379_),
    .B(_0720_),
    .Y(_1006_));
 sky130_fd_sc_hd__nand2_1 _4596_ (.A(_0384_),
    .B(_0350_),
    .Y(_1007_));
 sky130_fd_sc_hd__or2_1 _4597_ (.A(_0347_),
    .B(_0389_),
    .X(_1008_));
 sky130_fd_sc_hd__o2111a_1 _4598_ (.A1(_0711_),
    .A2(_0376_),
    .B1(_1006_),
    .C1(_1007_),
    .D1(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_1 _4599_ (.A(_0402_),
    .B(_0725_),
    .Y(_1010_));
 sky130_fd_sc_hd__nand2_1 _4600_ (.A(_0407_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1011_));
 sky130_fd_sc_hd__nand2_1 _4601_ (.A(_1010_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__a221oi_1 _4602_ (.A1(_0872_),
    .A2(_0395_),
    .B1(_0749_),
    .B2(_0399_),
    .C1(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__and4_1 _4603_ (.A(_1001_),
    .B(_1005_),
    .C(_1009_),
    .D(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__inv_2 _4604_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1015_));
 sky130_fd_sc_hd__o22ai_1 _4605_ (.A1(_0878_),
    .A2(_0423_),
    .B1(_1015_),
    .B2(_0426_),
    .Y(_1016_));
 sky130_fd_sc_hd__a221oi_1 _4606_ (.A1(_3110_),
    .A2(_0417_),
    .B1(_3113_),
    .B2(_0420_),
    .C1(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__nand2_1 _4607_ (.A(_0440_),
    .B(_3122_),
    .Y(_1018_));
 sky130_fd_sc_hd__o21ai_1 _4608_ (.A1(_0741_),
    .A2(_0437_),
    .B1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__a221oi_1 _4609_ (.A1(_3116_),
    .A2(_0431_),
    .B1(_3119_),
    .B2(_0434_),
    .C1(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__inv_2 _4610_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_1021_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_0455_),
    .B(_3093_),
    .Y(_1022_));
 sky130_fd_sc_hd__o21ai_1 _4612_ (.A1(_1021_),
    .A2(_0452_),
    .B1(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__a221oi_1 _4613_ (.A1(_3098_),
    .A2(_0446_),
    .B1(_3101_),
    .B2(_0449_),
    .C1(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__inv_2 _4614_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1025_));
 sky130_fd_sc_hd__o22ai_1 _4615_ (.A1(_0888_),
    .A2(_0467_),
    .B1(_1025_),
    .B2(_0470_),
    .Y(_1026_));
 sky130_fd_sc_hd__a221oi_1 _4616_ (.A1(_0787_),
    .A2(_0461_),
    .B1(_3284_),
    .B2(_0464_),
    .C1(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__and4_1 _4617_ (.A(_1017_),
    .B(_1020_),
    .C(_1024_),
    .D(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__o22ai_1 _4618_ (.A1(_0893_),
    .A2(_0487_),
    .B1(_0533_),
    .B2(_0490_),
    .Y(_1029_));
 sky130_fd_sc_hd__a221oi_1 _4619_ (.A1(_0892_),
    .A2(_0480_),
    .B1(_0525_),
    .B2(_0484_),
    .C1(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_0495_),
    .B(_0751_),
    .Y(_1031_));
 sky130_fd_sc_hd__buf_2 _4621_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_1032_));
 sky130_fd_sc_hd__nand2_1 _4622_ (.A(_0499_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _4623_ (.A(_0504_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1034_));
 sky130_fd_sc_hd__nand2_1 _4624_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_1035_));
 sky130_fd_sc_hd__and4_1 _4625_ (.A(_1031_),
    .B(_1033_),
    .C(_1034_),
    .D(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__o22ai_1 _4626_ (.A1(_0902_),
    .A2(_0513_),
    .B1(_0485_),
    .B2(_0516_),
    .Y(_1037_));
 sky130_fd_sc_hd__a22o_1 _4627_ (.A1(_0519_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .B1(_0521_),
    .B2(_0474_),
    .X(_1038_));
 sky130_fd_sc_hd__nor2_1 _4628_ (.A(_1037_),
    .B(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__inv_2 _4629_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_1040_));
 sky130_fd_sc_hd__o22ai_1 _4630_ (.A1(_0907_),
    .A2(_0535_),
    .B1(_1040_),
    .B2(_0538_),
    .Y(_1041_));
 sky130_fd_sc_hd__a221oi_1 _4631_ (.A1(_0569_),
    .A2(_0528_),
    .B1(_0580_),
    .B2(_0532_),
    .C1(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__and4_1 _4632_ (.A(_1030_),
    .B(_1036_),
    .C(_1039_),
    .D(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__nand2_1 _4633_ (.A(_0555_),
    .B(_0602_),
    .Y(_1044_));
 sky130_fd_sc_hd__nand2_1 _4634_ (.A(_0560_),
    .B(_0549_),
    .Y(_1045_));
 sky130_fd_sc_hd__nand2_1 _4635_ (.A(_1044_),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__a221oi_1 _4636_ (.A1(_0606_),
    .A2(_0548_),
    .B1(_0781_),
    .B2(_0552_),
    .C1(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__nand2_1 _4637_ (.A(_0574_),
    .B(_0595_),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_1 _4638_ (.A(_0579_),
    .B(_0774_),
    .Y(_1049_));
 sky130_fd_sc_hd__nand2_1 _4639_ (.A(_1048_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__a221oi_1 _4640_ (.A1(_0575_),
    .A2(_0568_),
    .B1(_0590_),
    .B2(_0571_),
    .C1(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__inv_2 _4641_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _4642_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_1053_));
 sky130_fd_sc_hd__nand2_1 _4643_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_1054_));
 sky130_fd_sc_hd__or2_1 _4644_ (.A(_0773_),
    .B(_0599_),
    .X(_1055_));
 sky130_fd_sc_hd__o2111a_1 _4645_ (.A1(_1052_),
    .A2(_0586_),
    .B1(_1053_),
    .C1(_1054_),
    .D1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_1 _4646_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_1057_));
 sky130_fd_sc_hd__o21ai_1 _4647_ (.A1(_0884_),
    .A2(_0612_),
    .B1(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__a221oi_2 _4648_ (.A1(_0924_),
    .A2(_0605_),
    .B1(_3072_),
    .B2(_0609_),
    .C1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__and4_1 _4649_ (.A(_1047_),
    .B(_1051_),
    .C(_1056_),
    .D(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__and4_1 _4650_ (.A(_1014_),
    .B(_1028_),
    .C(_1043_),
    .D(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__nand2_1 _4651_ (.A(_0624_),
    .B(_3291_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand3_1 _4652_ (.A(_0998_),
    .B(_1061_),
    .C(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__nor2_1 _4653_ (.A(_3134_),
    .B(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__nor2_1 _4654_ (.A(_0933_),
    .B(_1064_),
    .Y(_0294_));
 sky130_fd_sc_hd__o21ai_1 _4655_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_1065_));
 sky130_fd_sc_hd__inv_2 _4656_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_1066_));
 sky130_fd_sc_hd__nand2_1 _4657_ (.A(_3154_),
    .B(_3235_),
    .Y(_1067_));
 sky130_fd_sc_hd__a22o_1 _4658_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_1068_));
 sky130_fd_sc_hd__inv_2 _4659_ (.A(_1068_),
    .Y(_1069_));
 sky130_fd_sc_hd__o211a_1 _4660_ (.A1(_1066_),
    .A2(_3147_),
    .B1(_1067_),
    .C1(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__nand2_1 _4661_ (.A(_3190_),
    .B(_3195_),
    .Y(_1071_));
 sky130_fd_sc_hd__o21ai_1 _4662_ (.A1(_0642_),
    .A2(_3186_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__a221oi_1 _4663_ (.A1(_3212_),
    .A2(_3176_),
    .B1(_3214_),
    .B2(_3181_),
    .C1(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__nand2_1 _4664_ (.A(_3204_),
    .B(_0631_),
    .Y(_1074_));
 sky130_fd_sc_hd__nand2_1 _4665_ (.A(_3211_),
    .B(_3135_),
    .Y(_1075_));
 sky130_fd_sc_hd__or2_1 _4666_ (.A(_0630_),
    .B(_3219_),
    .X(_1076_));
 sky130_fd_sc_hd__o2111a_1 _4667_ (.A1(_0934_),
    .A2(_3200_),
    .B1(_1074_),
    .C1(_1075_),
    .D1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_1 _4668_ (.A(_3234_),
    .B(_3355_),
    .Y(_1078_));
 sky130_fd_sc_hd__nand2_1 _4669_ (.A(_3240_),
    .B(_3351_),
    .Y(_1079_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_1078_),
    .B(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__a221oi_1 _4671_ (.A1(_0675_),
    .A2(_3226_),
    .B1(_3365_),
    .B2(_3230_),
    .C1(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__and4_1 _4672_ (.A(_1070_),
    .B(_1073_),
    .C(_1077_),
    .D(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__nand2_1 _4673_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1083_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_3260_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_1084_));
 sky130_fd_sc_hd__or2_1 _4675_ (.A(_3268_),
    .B(_3265_),
    .X(_1085_));
 sky130_fd_sc_hd__o2111a_1 _4676_ (.A1(_3279_),
    .A2(_3252_),
    .B1(_1083_),
    .C1(_1084_),
    .D1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__nand2_1 _4677_ (.A(_3273_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1087_));
 sky130_fd_sc_hd__nand2_1 _4678_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1088_));
 sky130_fd_sc_hd__or2_1 _4679_ (.A(_3306_),
    .B(_3281_),
    .X(_1089_));
 sky130_fd_sc_hd__o2111a_1 _4680_ (.A1(_0820_),
    .A2(_3270_),
    .B1(_1087_),
    .C1(_1088_),
    .D1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__or2_1 _4681_ (.A(_3263_),
    .B(_3294_),
    .X(_1091_));
 sky130_fd_sc_hd__o221a_1 _4682_ (.A1(_0650_),
    .A2(_3287_),
    .B1(_3247_),
    .B2(_3290_),
    .C1(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__inv_2 _4683_ (.A(_3177_),
    .Y(_1093_));
 sky130_fd_sc_hd__o22ai_1 _4684_ (.A1(_0961_),
    .A2(_3305_),
    .B1(_1093_),
    .B2(_3308_),
    .Y(_1094_));
 sky130_fd_sc_hd__a221oi_1 _4685_ (.A1(_3182_),
    .A2(_3299_),
    .B1(_3191_),
    .B2(_3302_),
    .C1(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__and4_1 _4686_ (.A(_1086_),
    .B(_1090_),
    .C(_1092_),
    .D(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__inv_2 _4687_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_1097_));
 sky130_fd_sc_hd__o22ai_1 _4688_ (.A1(_0965_),
    .A2(_3324_),
    .B1(_1097_),
    .B2(_3328_),
    .Y(_1098_));
 sky130_fd_sc_hd__a221oi_1 _4689_ (.A1(_3331_),
    .A2(_3317_),
    .B1(_3335_),
    .B2(_3321_),
    .C1(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__nand2_1 _4690_ (.A(_3341_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _4691_ (.A(_3346_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2_1 _4692_ (.A(_1100_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__a221oi_1 _4693_ (.A1(_0681_),
    .A2(_3334_),
    .B1(_0834_),
    .B2(_3338_),
    .C1(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__nand2_1 _4694_ (.A(_3364_),
    .B(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_1104_));
 sky130_fd_sc_hd__o21ai_1 _4695_ (.A1(_0668_),
    .A2(_3361_),
    .B1(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__a221oi_1 _4696_ (.A1(_0677_),
    .A2(_3354_),
    .B1(_3325_),
    .B2(_3358_),
    .C1(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__buf_2 _4697_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_1107_));
 sky130_fd_sc_hd__nand2_1 _4698_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_1108_));
 sky130_fd_sc_hd__o21ai_1 _4699_ (.A1(_0990_),
    .A2(_3379_),
    .B1(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__a221oi_1 _4700_ (.A1(_0975_),
    .A2(_3372_),
    .B1(_1107_),
    .B2(_3376_),
    .C1(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__and4_1 _4701_ (.A(_1099_),
    .B(_1103_),
    .C(_1106_),
    .D(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__nand2_1 _4702_ (.A(_3393_),
    .B(_3416_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_1 _4703_ (.A(_3398_),
    .B(_0839_),
    .Y(_1113_));
 sky130_fd_sc_hd__or2_1 _4704_ (.A(_3406_),
    .B(_3403_),
    .X(_1114_));
 sky130_fd_sc_hd__o2111a_1 _4705_ (.A1(_3418_),
    .A2(_3390_),
    .B1(_1112_),
    .C1(_1113_),
    .D1(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__nand2_1 _4706_ (.A(_3411_),
    .B(_3440_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_3415_),
    .B(_0705_),
    .Y(_1117_));
 sky130_fd_sc_hd__or2_1 _4708_ (.A(_0844_),
    .B(_3420_),
    .X(_1118_));
 sky130_fd_sc_hd__o2111a_1 _4709_ (.A1(_0326_),
    .A2(_3408_),
    .B1(_1116_),
    .C1(_1117_),
    .D1(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__inv_2 _4710_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1120_));
 sky130_fd_sc_hd__nand2_1 _4711_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1121_));
 sky130_fd_sc_hd__o21ai_1 _4712_ (.A1(_1120_),
    .A2(_3433_),
    .B1(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__a221oi_1 _4713_ (.A1(_3394_),
    .A2(_3426_),
    .B1(_0687_),
    .B2(_3430_),
    .C1(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__nand2_1 _4714_ (.A(_0331_),
    .B(_0356_),
    .Y(_1124_));
 sky130_fd_sc_hd__o21ai_1 _4715_ (.A1(_1002_),
    .A2(_0328_),
    .B1(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__a221oi_1 _4716_ (.A1(_0854_),
    .A2(_3443_),
    .B1(_0370_),
    .B2(_0325_),
    .C1(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__and4_1 _4717_ (.A(_1115_),
    .B(_1119_),
    .C(_1123_),
    .D(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__and4_1 _4718_ (.A(_1082_),
    .B(_1096_),
    .C(_1111_),
    .D(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1129_));
 sky130_fd_sc_hd__o22ai_1 _4720_ (.A1(_0999_),
    .A2(_0349_),
    .B1(_1129_),
    .B2(_0353_),
    .Y(_1130_));
 sky130_fd_sc_hd__a221oi_1 _4721_ (.A1(_0392_),
    .A2(_0342_),
    .B1(_0396_),
    .B2(_0346_),
    .C1(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__inv_2 _4722_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(_0369_),
    .B(_0718_),
    .Y(_1133_));
 sky130_fd_sc_hd__o21ai_1 _4724_ (.A1(_1132_),
    .A2(_0366_),
    .B1(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__a221oi_1 _4725_ (.A1(_0385_),
    .A2(_0359_),
    .B1(_0720_),
    .B2(_0363_),
    .C1(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _4726_ (.A(_0379_),
    .B(_0868_),
    .Y(_1136_));
 sky130_fd_sc_hd__nand2_1 _4727_ (.A(_0384_),
    .B(_0337_),
    .Y(_1137_));
 sky130_fd_sc_hd__or2_1 _4728_ (.A(_0351_),
    .B(_0389_),
    .X(_1138_));
 sky130_fd_sc_hd__o2111a_1 _4729_ (.A1(_0860_),
    .A2(_0376_),
    .B1(_1136_),
    .C1(_1137_),
    .D1(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(_0402_),
    .B(_0872_),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(_0407_),
    .B(_0725_),
    .Y(_1141_));
 sky130_fd_sc_hd__nand2_1 _4732_ (.A(_1140_),
    .B(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__a221oi_1 _4733_ (.A1(_0749_),
    .A2(_0395_),
    .B1(_0500_),
    .B2(_0399_),
    .C1(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__and4_1 _4734_ (.A(_1131_),
    .B(_1135_),
    .C(_1139_),
    .D(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__inv_2 _4735_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1145_));
 sky130_fd_sc_hd__o22ai_1 _4736_ (.A1(_1015_),
    .A2(_0423_),
    .B1(_1145_),
    .B2(_0426_),
    .Y(_1146_));
 sky130_fd_sc_hd__a221oi_1 _4737_ (.A1(_3113_),
    .A2(_0417_),
    .B1(_3116_),
    .B2(_0420_),
    .C1(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0440_),
    .B(_3125_),
    .Y(_1148_));
 sky130_fd_sc_hd__o21ai_1 _4739_ (.A1(_0888_),
    .A2(_0437_),
    .B1(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__a221oi_1 _4740_ (.A1(_3119_),
    .A2(_0431_),
    .B1(_3122_),
    .B2(_0434_),
    .C1(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_1 _4741_ (.A(_0455_),
    .B(_3098_),
    .Y(_1151_));
 sky130_fd_sc_hd__o21ai_1 _4742_ (.A1(_0421_),
    .A2(_0452_),
    .B1(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__a221oi_1 _4743_ (.A1(_3101_),
    .A2(_0446_),
    .B1(_3104_),
    .B2(_0449_),
    .C1(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__o22ai_1 _4744_ (.A1(_1025_),
    .A2(_0467_),
    .B1(_3288_),
    .B2(_0470_),
    .Y(_1154_));
 sky130_fd_sc_hd__a221oi_1 _4745_ (.A1(_3284_),
    .A2(_0461_),
    .B1(_3291_),
    .B2(_0464_),
    .C1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__and4_1 _4746_ (.A(_1147_),
    .B(_1150_),
    .C(_1153_),
    .D(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__o22ai_1 _4747_ (.A1(_0533_),
    .A2(_0487_),
    .B1(_0536_),
    .B2(_0490_),
    .Y(_1157_));
 sky130_fd_sc_hd__a221oi_1 _4748_ (.A1(_0525_),
    .A2(_0480_),
    .B1(_0529_),
    .B2(_0484_),
    .C1(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__nand2_1 _4749_ (.A(_0495_),
    .B(_0897_),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_1 _4750_ (.A(_0499_),
    .B(_0522_),
    .Y(_1160_));
 sky130_fd_sc_hd__nand2_1 _4751_ (.A(_0504_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_1162_));
 sky130_fd_sc_hd__and4_1 _4753_ (.A(_1159_),
    .B(_1160_),
    .C(_1161_),
    .D(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__o22ai_1 _4754_ (.A1(_0485_),
    .A2(_0513_),
    .B1(_0488_),
    .B2(_0516_),
    .Y(_1164_));
 sky130_fd_sc_hd__a22o_1 _4755_ (.A1(_0519_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .B1(_0521_),
    .B2(_0481_),
    .X(_1165_));
 sky130_fd_sc_hd__nor2_1 _4756_ (.A(_1164_),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__inv_2 _4757_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_1167_));
 sky130_fd_sc_hd__o22ai_1 _4758_ (.A1(_1040_),
    .A2(_0535_),
    .B1(_1167_),
    .B2(_0538_),
    .Y(_1168_));
 sky130_fd_sc_hd__a221oi_1 _4759_ (.A1(_0580_),
    .A2(_0528_),
    .B1(_0575_),
    .B2(_0532_),
    .C1(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__and4_1 _4760_ (.A(_1158_),
    .B(_1163_),
    .C(_1166_),
    .D(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nand2_1 _4761_ (.A(_0555_),
    .B(_0606_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(_0560_),
    .B(_0602_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _4763_ (.A(_1171_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__a221oi_1 _4764_ (.A1(_0781_),
    .A2(_0548_),
    .B1(_0924_),
    .B2(_0552_),
    .C1(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_1 _4765_ (.A(_0574_),
    .B(_0776_),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _4766_ (.A(_0579_),
    .B(_0595_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _4767_ (.A(_1175_),
    .B(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__a221oi_1 _4768_ (.A1(_0590_),
    .A2(_0568_),
    .B1(_0774_),
    .B2(_0571_),
    .C1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__inv_2 _4769_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1179_));
 sky130_fd_sc_hd__nand2_1 _4770_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_1180_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1181_));
 sky130_fd_sc_hd__or2_1 _4772_ (.A(_0919_),
    .B(_0599_),
    .X(_1182_));
 sky130_fd_sc_hd__o2111a_1 _4773_ (.A1(_1179_),
    .A2(_0586_),
    .B1(_1180_),
    .C1(_1181_),
    .D1(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_1184_));
 sky130_fd_sc_hd__o21ai_1 _4775_ (.A1(_1021_),
    .A2(_0612_),
    .B1(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__a221oi_1 _4776_ (.A1(_3072_),
    .A2(_0605_),
    .B1(_3084_),
    .B2(_0609_),
    .C1(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__and4_1 _4777_ (.A(_1174_),
    .B(_1178_),
    .C(_1183_),
    .D(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__and4_1 _4778_ (.A(_1144_),
    .B(_1156_),
    .C(_1170_),
    .D(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(_0624_),
    .B(_3261_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand3_1 _4780_ (.A(_1128_),
    .B(_1188_),
    .C(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_1 _4781_ (.A(_3134_),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__nor2_1 _4782_ (.A(_1065_),
    .B(_1191_),
    .Y(_0293_));
 sky130_fd_sc_hd__o21ai_1 _4783_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_1192_));
 sky130_fd_sc_hd__inv_2 _4784_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_1193_));
 sky130_fd_sc_hd__nand2_1 _4785_ (.A(_3154_),
    .B(_3222_),
    .Y(_1194_));
 sky130_fd_sc_hd__a22o_1 _4786_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_1195_));
 sky130_fd_sc_hd__inv_2 _4787_ (.A(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__o211a_1 _4788_ (.A1(_1193_),
    .A2(_3147_),
    .B1(_1194_),
    .C1(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_3190_),
    .B(_3135_),
    .Y(_1198_));
 sky130_fd_sc_hd__o21ai_1 _4790_ (.A1(_3196_),
    .A2(_3186_),
    .B1(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__a221oi_1 _4791_ (.A1(_3214_),
    .A2(_3176_),
    .B1(_3205_),
    .B2(_3181_),
    .C1(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nand2_1 _4792_ (.A(_3204_),
    .B(_3167_),
    .Y(_1201_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_3211_),
    .B(_3155_),
    .Y(_1202_));
 sky130_fd_sc_hd__or2_1 _4794_ (.A(_0792_),
    .B(_3219_),
    .X(_1203_));
 sky130_fd_sc_hd__o2111a_1 _4795_ (.A1(_1066_),
    .A2(_3200_),
    .B1(_1201_),
    .C1(_1202_),
    .D1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__nand2_1 _4796_ (.A(_3234_),
    .B(_0675_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(_3240_),
    .B(_3355_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand2_1 _4798_ (.A(_1205_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__a221oi_1 _4799_ (.A1(_3365_),
    .A2(_3226_),
    .B1(_0677_),
    .B2(_3230_),
    .C1(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__and4_1 _4800_ (.A(_1197_),
    .B(_1200_),
    .C(_1204_),
    .D(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__nand2_1 _4801_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1210_));
 sky130_fd_sc_hd__nand2_1 _4802_ (.A(_3260_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1211_));
 sky130_fd_sc_hd__or2_1 _4803_ (.A(_3303_),
    .B(_3265_),
    .X(_1212_));
 sky130_fd_sc_hd__o2111a_1 _4804_ (.A1(_0658_),
    .A2(_3252_),
    .B1(_1210_),
    .C1(_1211_),
    .D1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__nand2_1 _4805_ (.A(_3273_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _4806_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1215_));
 sky130_fd_sc_hd__or2_1 _4807_ (.A(_0664_),
    .B(_3281_),
    .X(_1216_));
 sky130_fd_sc_hd__o2111a_1 _4808_ (.A1(_0961_),
    .A2(_3270_),
    .B1(_1214_),
    .C1(_1215_),
    .D1(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__or2_1 _4809_ (.A(_0653_),
    .B(_3294_),
    .X(_1218_));
 sky130_fd_sc_hd__o221a_1 _4810_ (.A1(_3263_),
    .A2(_3287_),
    .B1(_0650_),
    .B2(_3290_),
    .C1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__o22ai_1 _4811_ (.A1(_1093_),
    .A2(_3305_),
    .B1(_3183_),
    .B2(_3308_),
    .Y(_1220_));
 sky130_fd_sc_hd__a221oi_1 _4812_ (.A1(_3191_),
    .A2(_3299_),
    .B1(_3212_),
    .B2(_3302_),
    .C1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__and4_1 _4813_ (.A(_1213_),
    .B(_1217_),
    .C(_1219_),
    .D(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__inv_2 _4814_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1223_));
 sky130_fd_sc_hd__o22ai_1 _4815_ (.A1(_1097_),
    .A2(_3324_),
    .B1(_1223_),
    .B2(_3328_),
    .Y(_1224_));
 sky130_fd_sc_hd__a221oi_1 _4816_ (.A1(_3335_),
    .A2(_3317_),
    .B1(_3369_),
    .B2(_3321_),
    .C1(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__nand2_1 _4817_ (.A(_3341_),
    .B(_0681_),
    .Y(_1226_));
 sky130_fd_sc_hd__nand2_1 _4818_ (.A(_3346_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1227_));
 sky130_fd_sc_hd__nand2_1 _4819_ (.A(_1226_),
    .B(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__a221oi_1 _4820_ (.A1(_0834_),
    .A2(_3334_),
    .B1(_0975_),
    .B2(_3338_),
    .C1(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(_3364_),
    .B(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_1230_));
 sky130_fd_sc_hd__o21ai_1 _4822_ (.A1(_0824_),
    .A2(_3361_),
    .B1(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__a221oi_1 _4823_ (.A1(_3325_),
    .A2(_3354_),
    .B1(_3312_),
    .B2(_3358_),
    .C1(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2_1 _4824_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_1233_));
 sky130_fd_sc_hd__o21ai_1 _4825_ (.A1(_1120_),
    .A2(_3379_),
    .B1(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__a221oi_1 _4826_ (.A1(_1107_),
    .A2(_3372_),
    .B1(_3423_),
    .B2(_3376_),
    .C1(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__and4_1 _4827_ (.A(_1225_),
    .B(_1229_),
    .C(_1232_),
    .D(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__nand2_1 _4828_ (.A(_3393_),
    .B(_0696_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _4829_ (.A(_3398_),
    .B(_0980_),
    .Y(_1238_));
 sky130_fd_sc_hd__or2_1 _4830_ (.A(_0694_),
    .B(_3403_),
    .X(_1239_));
 sky130_fd_sc_hd__o2111a_1 _4831_ (.A1(_0698_),
    .A2(_3390_),
    .B1(_1237_),
    .C1(_1238_),
    .D1(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_3411_),
    .B(_0322_),
    .Y(_1241_));
 sky130_fd_sc_hd__nand2_1 _4833_ (.A(_3415_),
    .B(_0853_),
    .Y(_1242_));
 sky130_fd_sc_hd__or2_1 _4834_ (.A(_0985_),
    .B(_3420_),
    .X(_1243_));
 sky130_fd_sc_hd__o2111a_1 _4835_ (.A1(_0364_),
    .A2(_3408_),
    .B1(_1241_),
    .C1(_1242_),
    .D1(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__nand2_1 _4836_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1245_));
 sky130_fd_sc_hd__o21ai_1 _4837_ (.A1(_3387_),
    .A2(_3433_),
    .B1(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a221oi_1 _4838_ (.A1(_0687_),
    .A2(_3426_),
    .B1(_0839_),
    .B2(_3430_),
    .C1(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_0331_),
    .B(_0360_),
    .Y(_1248_));
 sky130_fd_sc_hd__o21ai_1 _4840_ (.A1(_1132_),
    .A2(_0328_),
    .B1(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__a221oi_1 _4841_ (.A1(_0370_),
    .A2(_3443_),
    .B1(_0356_),
    .B2(_0325_),
    .C1(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__and4_1 _4842_ (.A(_1240_),
    .B(_1244_),
    .C(_1247_),
    .D(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__and4_1 _4843_ (.A(_1209_),
    .B(_1222_),
    .C(_1236_),
    .D(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__inv_2 _4844_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1253_));
 sky130_fd_sc_hd__o22ai_1 _4845_ (.A1(_1129_),
    .A2(_0349_),
    .B1(_1253_),
    .B2(_0353_),
    .Y(_1254_));
 sky130_fd_sc_hd__a221oi_1 _4846_ (.A1(_0396_),
    .A2(_0342_),
    .B1(_0725_),
    .B2(_0346_),
    .C1(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(_0369_),
    .B(_0385_),
    .Y(_1256_));
 sky130_fd_sc_hd__o21ai_1 _4848_ (.A1(_0387_),
    .A2(_0366_),
    .B1(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__a221oi_1 _4849_ (.A1(_0720_),
    .A2(_0359_),
    .B1(_0868_),
    .B2(_0363_),
    .C1(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_0379_),
    .B(_0350_),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_1 _4851_ (.A(_0384_),
    .B(_0343_),
    .Y(_1260_));
 sky130_fd_sc_hd__or2_1 _4852_ (.A(_0711_),
    .B(_0389_),
    .X(_1261_));
 sky130_fd_sc_hd__o2111a_1 _4853_ (.A1(_0999_),
    .A2(_0376_),
    .B1(_1259_),
    .C1(_1260_),
    .D1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_0402_),
    .B(_0749_),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_0407_),
    .B(_0872_),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_1 _4856_ (.A(_1263_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__a221oi_1 _4857_ (.A1(_0500_),
    .A2(_0395_),
    .B1(_0751_),
    .B2(_0399_),
    .C1(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__and4_1 _4858_ (.A(_1255_),
    .B(_1258_),
    .C(_1262_),
    .D(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__inv_2 _4859_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1268_));
 sky130_fd_sc_hd__o22ai_1 _4860_ (.A1(_1145_),
    .A2(_0423_),
    .B1(_1268_),
    .B2(_0426_),
    .Y(_1269_));
 sky130_fd_sc_hd__a221oi_1 _4861_ (.A1(_3116_),
    .A2(_0417_),
    .B1(_3119_),
    .B2(_0420_),
    .C1(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__nand2_1 _4862_ (.A(_0440_),
    .B(_3129_),
    .Y(_1271_));
 sky130_fd_sc_hd__o21ai_1 _4863_ (.A1(_1025_),
    .A2(_0437_),
    .B1(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__a221oi_1 _4864_ (.A1(_3122_),
    .A2(_0431_),
    .B1(_3125_),
    .B2(_0434_),
    .C1(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1274_));
 sky130_fd_sc_hd__o21ai_1 _4866_ (.A1(_0424_),
    .A2(_0452_),
    .B1(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__a221oi_1 _4867_ (.A1(_3104_),
    .A2(_0446_),
    .B1(_3107_),
    .B2(_0449_),
    .C1(_1275_),
    .Y(_1276_));
 sky130_fd_sc_hd__o22ai_1 _4868_ (.A1(_3288_),
    .A2(_0467_),
    .B1(_3285_),
    .B2(_0470_),
    .Y(_1277_));
 sky130_fd_sc_hd__a221oi_1 _4869_ (.A1(_3291_),
    .A2(_0461_),
    .B1(_3261_),
    .B2(_0464_),
    .C1(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__and4_1 _4870_ (.A(_1270_),
    .B(_1273_),
    .C(_1276_),
    .D(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__o22ai_1 _4871_ (.A1(_0536_),
    .A2(_0487_),
    .B1(_0761_),
    .B2(_0490_),
    .Y(_1280_));
 sky130_fd_sc_hd__a221oi_1 _4872_ (.A1(_0529_),
    .A2(_0480_),
    .B1(_0565_),
    .B2(_0484_),
    .C1(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_0495_),
    .B(_1032_),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2_1 _4874_ (.A(_0499_),
    .B(_0758_),
    .Y(_1283_));
 sky130_fd_sc_hd__nand2_1 _4875_ (.A(_0504_),
    .B(_0897_),
    .Y(_1284_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1285_));
 sky130_fd_sc_hd__and4_1 _4877_ (.A(_1282_),
    .B(_1283_),
    .C(_1284_),
    .D(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__o22ai_1 _4878_ (.A1(_0488_),
    .A2(_0513_),
    .B1(_0746_),
    .B2(_0516_),
    .Y(_1287_));
 sky130_fd_sc_hd__a22o_1 _4879_ (.A1(_0519_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .B1(_0521_),
    .B2(_0745_),
    .X(_1288_));
 sky130_fd_sc_hd__nor2_1 _4880_ (.A(_1287_),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__inv_2 _4881_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .Y(_1290_));
 sky130_fd_sc_hd__o22ai_1 _4882_ (.A1(_1167_),
    .A2(_0535_),
    .B1(_1290_),
    .B2(_0538_),
    .Y(_1291_));
 sky130_fd_sc_hd__a221oi_1 _4883_ (.A1(_0575_),
    .A2(_0528_),
    .B1(_0590_),
    .B2(_0532_),
    .C1(_1291_),
    .Y(_1292_));
 sky130_fd_sc_hd__and4_1 _4884_ (.A(_1281_),
    .B(_1286_),
    .C(_1289_),
    .D(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(_0555_),
    .B(_0781_),
    .Y(_1294_));
 sky130_fd_sc_hd__nand2_1 _4886_ (.A(_0560_),
    .B(_0606_),
    .Y(_1295_));
 sky130_fd_sc_hd__nand2_1 _4887_ (.A(_1294_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__a221oi_1 _4888_ (.A1(_0924_),
    .A2(_0548_),
    .B1(_3072_),
    .B2(_0552_),
    .C1(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__nand2_1 _4889_ (.A(_0574_),
    .B(_0561_),
    .Y(_1298_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(_0579_),
    .B(_0776_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_1298_),
    .B(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__a221oi_2 _4892_ (.A1(_0774_),
    .A2(_0568_),
    .B1(_0595_),
    .B2(_0571_),
    .C1(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_2 _4893_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1302_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_1303_));
 sky130_fd_sc_hd__nand2_1 _4895_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1304_));
 sky130_fd_sc_hd__or2_1 _4896_ (.A(_1052_),
    .B(_0599_),
    .X(_1305_));
 sky130_fd_sc_hd__o2111a_1 _4897_ (.A1(_1302_),
    .A2(_0586_),
    .B1(_1303_),
    .C1(_1304_),
    .D1(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_1307_));
 sky130_fd_sc_hd__o21ai_1 _4899_ (.A1(_0421_),
    .A2(_0612_),
    .B1(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__a221oi_1 _4900_ (.A1(_3084_),
    .A2(_0605_),
    .B1(_3087_),
    .B2(_0609_),
    .C1(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__and4_1 _4901_ (.A(_1297_),
    .B(_1301_),
    .C(_1306_),
    .D(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__and4_1 _4902_ (.A(_1267_),
    .B(_1279_),
    .C(_1293_),
    .D(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__nand2_1 _4903_ (.A(_0624_),
    .B(_3246_),
    .Y(_1312_));
 sky130_fd_sc_hd__nand3_1 _4904_ (.A(_1252_),
    .B(_1311_),
    .C(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__nor2_1 _4905_ (.A(_3134_),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__nor2_1 _4906_ (.A(_1192_),
    .B(_1314_),
    .Y(_0292_));
 sky130_fd_sc_hd__o21ai_1 _4907_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_1315_));
 sky130_fd_sc_hd__inv_2 _4908_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2_1 _4909_ (.A(_3154_),
    .B(_3227_),
    .Y(_1317_));
 sky130_fd_sc_hd__a22o_1 _4910_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_1318_));
 sky130_fd_sc_hd__inv_2 _4911_ (.A(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__o211a_1 _4912_ (.A1(_1316_),
    .A2(_3147_),
    .B1(_1317_),
    .C1(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__nand2_1 _4913_ (.A(_3190_),
    .B(_3155_),
    .Y(_1321_));
 sky130_fd_sc_hd__o21ai_1 _4914_ (.A1(_3136_),
    .A2(_3186_),
    .B1(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__a221oi_1 _4915_ (.A1(_3205_),
    .A2(_3176_),
    .B1(_3195_),
    .B2(_3181_),
    .C1(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(_3204_),
    .B(_3241_),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _4917_ (.A(_3211_),
    .B(_0631_),
    .Y(_1325_));
 sky130_fd_sc_hd__or2_1 _4918_ (.A(_0934_),
    .B(_3219_),
    .X(_1326_));
 sky130_fd_sc_hd__o2111a_1 _4919_ (.A1(_1193_),
    .A2(_3200_),
    .B1(_1324_),
    .C1(_1325_),
    .D1(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__nand2_1 _4920_ (.A(_3234_),
    .B(_3365_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2_1 _4921_ (.A(_3240_),
    .B(_0675_),
    .Y(_1329_));
 sky130_fd_sc_hd__nand2_1 _4922_ (.A(_1328_),
    .B(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__a221oi_1 _4923_ (.A1(_0677_),
    .A2(_3226_),
    .B1(_3325_),
    .B2(_3230_),
    .C1(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__and4_1 _4924_ (.A(_1320_),
    .B(_1323_),
    .C(_1327_),
    .D(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__nand2_1 _4925_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_1 _4926_ (.A(_3260_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1334_));
 sky130_fd_sc_hd__or2_1 _4927_ (.A(_3306_),
    .B(_3265_),
    .X(_1335_));
 sky130_fd_sc_hd__o2111a_1 _4928_ (.A1(_3268_),
    .A2(_3252_),
    .B1(_1333_),
    .C1(_1334_),
    .D1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__nand2_1 _4929_ (.A(_3273_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1338_));
 sky130_fd_sc_hd__or2_1 _4931_ (.A(_0820_),
    .B(_3281_),
    .X(_1339_));
 sky130_fd_sc_hd__o2111a_1 _4932_ (.A1(_1093_),
    .A2(_3270_),
    .B1(_1337_),
    .C1(_1338_),
    .D1(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__or2_1 _4933_ (.A(_3279_),
    .B(_3294_),
    .X(_1341_));
 sky130_fd_sc_hd__o221a_1 _4934_ (.A1(_0653_),
    .A2(_3287_),
    .B1(_3263_),
    .B2(_3290_),
    .C1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__o22ai_1 _4935_ (.A1(_3183_),
    .A2(_3305_),
    .B1(_0636_),
    .B2(_3308_),
    .Y(_1343_));
 sky130_fd_sc_hd__a221oi_1 _4936_ (.A1(_3212_),
    .A2(_3299_),
    .B1(_3214_),
    .B2(_3302_),
    .C1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__and4_1 _4937_ (.A(_1336_),
    .B(_1340_),
    .C(_1342_),
    .D(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__inv_2 _4938_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_1346_));
 sky130_fd_sc_hd__o22ai_1 _4939_ (.A1(_1223_),
    .A2(_3324_),
    .B1(_1346_),
    .B2(_3328_),
    .Y(_1347_));
 sky130_fd_sc_hd__a221oi_1 _4940_ (.A1(_3369_),
    .A2(_3317_),
    .B1(_3373_),
    .B2(_3321_),
    .C1(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__nand2_1 _4941_ (.A(_3341_),
    .B(_0834_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(_3346_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4943_ (.A(_1349_),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__a221oi_1 _4944_ (.A1(_0975_),
    .A2(_3334_),
    .B1(_1107_),
    .B2(_3338_),
    .C1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__nand2_1 _4945_ (.A(_3364_),
    .B(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_1353_));
 sky130_fd_sc_hd__o21ai_1 _4946_ (.A1(_0965_),
    .A2(_3361_),
    .B1(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__a221oi_1 _4947_ (.A1(_3312_),
    .A2(_3354_),
    .B1(_3318_),
    .B2(_3358_),
    .C1(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_1 _4948_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1356_));
 sky130_fd_sc_hd__o21ai_1 _4949_ (.A1(_3387_),
    .A2(_3379_),
    .B1(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__a221oi_1 _4950_ (.A1(_3423_),
    .A2(_3372_),
    .B1(_3427_),
    .B2(_3376_),
    .C1(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__and4_1 _4951_ (.A(_1348_),
    .B(_1352_),
    .C(_1355_),
    .D(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__nand2_1 _4952_ (.A(_3393_),
    .B(_3440_),
    .Y(_1360_));
 sky130_fd_sc_hd__nand2_1 _4953_ (.A(_3398_),
    .B(_3416_),
    .Y(_1361_));
 sky130_fd_sc_hd__or2_1 _4954_ (.A(_0844_),
    .B(_3403_),
    .X(_1362_));
 sky130_fd_sc_hd__o2111a_1 _4955_ (.A1(_3406_),
    .A2(_3390_),
    .B1(_1360_),
    .C1(_1361_),
    .D1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__nand2_1 _4956_ (.A(_3411_),
    .B(_0705_),
    .Y(_1364_));
 sky130_fd_sc_hd__nand2_1 _4957_ (.A(_3415_),
    .B(_0854_),
    .Y(_1365_));
 sky130_fd_sc_hd__or2_1 _4958_ (.A(_0326_),
    .B(_3420_),
    .X(_1366_));
 sky130_fd_sc_hd__o2111a_1 _4959_ (.A1(_0714_),
    .A2(_3408_),
    .B1(_1364_),
    .C1(_1365_),
    .D1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__nand2_1 _4960_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1368_));
 sky130_fd_sc_hd__o21ai_1 _4961_ (.A1(_0686_),
    .A2(_3433_),
    .B1(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__a221oi_1 _4962_ (.A1(_0839_),
    .A2(_3426_),
    .B1(_0980_),
    .B2(_3430_),
    .C1(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__nand2_1 _4963_ (.A(_0331_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1371_));
 sky130_fd_sc_hd__o21ai_1 _4964_ (.A1(_0387_),
    .A2(_0328_),
    .B1(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__a221oi_1 _4965_ (.A1(_0356_),
    .A2(_3443_),
    .B1(_0360_),
    .B2(_0325_),
    .C1(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__and4_1 _4966_ (.A(_1363_),
    .B(_1367_),
    .C(_1370_),
    .D(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__and4_1 _4967_ (.A(_1332_),
    .B(_1345_),
    .C(_1359_),
    .D(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__inv_2 _4968_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1376_));
 sky130_fd_sc_hd__o22ai_1 _4969_ (.A1(_1253_),
    .A2(_0349_),
    .B1(_1376_),
    .B2(_0353_),
    .Y(_1377_));
 sky130_fd_sc_hd__a221oi_1 _4970_ (.A1(_0725_),
    .A2(_0342_),
    .B1(_0872_),
    .B2(_0346_),
    .C1(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_0369_),
    .B(_0720_),
    .Y(_1379_));
 sky130_fd_sc_hd__o21ai_1 _4972_ (.A1(_0722_),
    .A2(_0366_),
    .B1(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__a221oi_1 _4973_ (.A1(_0868_),
    .A2(_0359_),
    .B1(_0350_),
    .B2(_0363_),
    .C1(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_0379_),
    .B(_0337_),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _4975_ (.A(_0384_),
    .B(_0408_),
    .Y(_1383_));
 sky130_fd_sc_hd__or2_1 _4976_ (.A(_0860_),
    .B(_0389_),
    .X(_1384_));
 sky130_fd_sc_hd__o2111a_1 _4977_ (.A1(_1129_),
    .A2(_0376_),
    .B1(_1382_),
    .C1(_1383_),
    .D1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(_0402_),
    .B(_0500_),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_0407_),
    .B(_0749_),
    .Y(_1387_));
 sky130_fd_sc_hd__nand2_1 _4980_ (.A(_1386_),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__a221oi_1 _4981_ (.A1(_0751_),
    .A2(_0395_),
    .B1(_0897_),
    .B2(_0399_),
    .C1(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__and4_1 _4982_ (.A(_1378_),
    .B(_1381_),
    .C(_1385_),
    .D(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__o22ai_1 _4983_ (.A1(_1268_),
    .A2(_0423_),
    .B1(_0435_),
    .B2(_0426_),
    .Y(_1391_));
 sky130_fd_sc_hd__a221oi_1 _4984_ (.A1(_3119_),
    .A2(_0417_),
    .B1(_3122_),
    .B2(_0420_),
    .C1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__nand2_1 _4985_ (.A(_0440_),
    .B(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1393_));
 sky130_fd_sc_hd__o21ai_1 _4986_ (.A1(_3288_),
    .A2(_0437_),
    .B1(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__a221oi_1 _4987_ (.A1(_3125_),
    .A2(_0431_),
    .B1(_3129_),
    .B2(_0434_),
    .C1(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_1396_));
 sky130_fd_sc_hd__o21ai_1 _4989_ (.A1(_0731_),
    .A2(_0452_),
    .B1(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__a221oi_1 _4990_ (.A1(_3107_),
    .A2(_0446_),
    .B1(_3110_),
    .B2(_0449_),
    .C1(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__o22ai_1 _4991_ (.A1(_3285_),
    .A2(_0467_),
    .B1(_3292_),
    .B2(_0470_),
    .Y(_1399_));
 sky130_fd_sc_hd__a221oi_1 _4992_ (.A1(_3261_),
    .A2(_0461_),
    .B1(_3246_),
    .B2(_0464_),
    .C1(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__and4_1 _4993_ (.A(_1392_),
    .B(_1395_),
    .C(_1398_),
    .D(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__o22ai_1 _4994_ (.A1(_0761_),
    .A2(_0487_),
    .B1(_0907_),
    .B2(_0490_),
    .Y(_1402_));
 sky130_fd_sc_hd__a221oi_1 _4995_ (.A1(_0565_),
    .A2(_0480_),
    .B1(_0569_),
    .B2(_0484_),
    .C1(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__nand2_1 _4996_ (.A(_0495_),
    .B(_0522_),
    .Y(_1404_));
 sky130_fd_sc_hd__nand2_1 _4997_ (.A(_0499_),
    .B(_0904_),
    .Y(_1405_));
 sky130_fd_sc_hd__nand2_1 _4998_ (.A(_0504_),
    .B(_1032_),
    .Y(_1406_));
 sky130_fd_sc_hd__nand2_1 _4999_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1407_));
 sky130_fd_sc_hd__and4_1 _5000_ (.A(_1404_),
    .B(_1405_),
    .C(_1406_),
    .D(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__o22ai_1 _5001_ (.A1(_0746_),
    .A2(_0513_),
    .B1(_0893_),
    .B2(_0516_),
    .Y(_1409_));
 sky130_fd_sc_hd__a22o_1 _5002_ (.A1(_0519_),
    .A2(_0745_),
    .B1(_0521_),
    .B2(_0892_),
    .X(_1410_));
 sky130_fd_sc_hd__nor2_1 _5003_ (.A(_1409_),
    .B(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__inv_2 _5004_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .Y(_1412_));
 sky130_fd_sc_hd__o22ai_1 _5005_ (.A1(_1290_),
    .A2(_0535_),
    .B1(_1412_),
    .B2(_0538_),
    .Y(_1413_));
 sky130_fd_sc_hd__a221oi_1 _5006_ (.A1(_0590_),
    .A2(_0528_),
    .B1(_0774_),
    .B2(_0532_),
    .C1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__and4_1 _5007_ (.A(_1403_),
    .B(_1408_),
    .C(_1411_),
    .D(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_0555_),
    .B(_0924_),
    .Y(_1416_));
 sky130_fd_sc_hd__nand2_1 _5009_ (.A(_0560_),
    .B(_0781_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(_1416_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__a221oi_1 _5011_ (.A1(_3072_),
    .A2(_0548_),
    .B1(_3084_),
    .B2(_0552_),
    .C1(_1418_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _5012_ (.A(_0574_),
    .B(_0556_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _5013_ (.A(_0579_),
    .B(_0561_),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _5014_ (.A(_1420_),
    .B(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__a221oi_1 _5015_ (.A1(_0595_),
    .A2(_0568_),
    .B1(_0776_),
    .B2(_0571_),
    .C1(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__inv_2 _5016_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1424_));
 sky130_fd_sc_hd__nand2_1 _5017_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1425_));
 sky130_fd_sc_hd__nand2_1 _5018_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1426_));
 sky130_fd_sc_hd__or2_1 _5019_ (.A(_1179_),
    .B(_0599_),
    .X(_1427_));
 sky130_fd_sc_hd__o2111a_1 _5020_ (.A1(_1424_),
    .A2(_0586_),
    .B1(_1425_),
    .C1(_1426_),
    .D1(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__nand2_1 _5021_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_1429_));
 sky130_fd_sc_hd__o21ai_1 _5022_ (.A1(_0424_),
    .A2(_0612_),
    .B1(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__a221oi_1 _5023_ (.A1(_3087_),
    .A2(_0605_),
    .B1(_3090_),
    .B2(_0609_),
    .C1(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__and4_1 _5024_ (.A(_1419_),
    .B(_1423_),
    .C(_1428_),
    .D(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__and4_1 _5025_ (.A(_1390_),
    .B(_1401_),
    .C(_1415_),
    .D(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_0624_),
    .B(_3256_),
    .Y(_1434_));
 sky130_fd_sc_hd__nand3_1 _5027_ (.A(_1375_),
    .B(_1433_),
    .C(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__nor2_1 _5028_ (.A(_3134_),
    .B(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hd__nor2_1 _5029_ (.A(_1315_),
    .B(_1436_),
    .Y(_0291_));
 sky130_fd_sc_hd__o21ai_1 _5030_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_1437_));
 sky130_fd_sc_hd__inv_2 _5031_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .Y(_1438_));
 sky130_fd_sc_hd__nand2_1 _5032_ (.A(_3154_),
    .B(_3351_),
    .Y(_1439_));
 sky130_fd_sc_hd__a22o_1 _5033_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_1440_));
 sky130_fd_sc_hd__inv_2 _5034_ (.A(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__o211a_1 _5035_ (.A1(_1438_),
    .A2(_3147_),
    .B1(_1439_),
    .C1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__nand2_1 _5036_ (.A(_3190_),
    .B(_0631_),
    .Y(_1443_));
 sky130_fd_sc_hd__o21ai_1 _5037_ (.A1(_0630_),
    .A2(_3186_),
    .B1(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__a221oi_1 _5038_ (.A1(_3195_),
    .A2(_3176_),
    .B1(_3135_),
    .B2(_3181_),
    .C1(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(_3204_),
    .B(_3235_),
    .Y(_1446_));
 sky130_fd_sc_hd__nand2_1 _5040_ (.A(_3211_),
    .B(_3167_),
    .Y(_1447_));
 sky130_fd_sc_hd__or2_1 _5041_ (.A(_1066_),
    .B(_3219_),
    .X(_1448_));
 sky130_fd_sc_hd__o2111a_1 _5042_ (.A1(_1316_),
    .A2(_3200_),
    .B1(_1446_),
    .C1(_1447_),
    .D1(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__nand2_1 _5043_ (.A(_3234_),
    .B(_0677_),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _5044_ (.A(_3240_),
    .B(_3365_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_1 _5045_ (.A(_1450_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__a221oi_1 _5046_ (.A1(_3325_),
    .A2(_3226_),
    .B1(_3312_),
    .B2(_3230_),
    .C1(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__and4_1 _5047_ (.A(_1442_),
    .B(_1445_),
    .C(_1449_),
    .D(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1455_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_3260_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1456_));
 sky130_fd_sc_hd__or2_1 _5050_ (.A(_0664_),
    .B(_3265_),
    .X(_1457_));
 sky130_fd_sc_hd__o2111a_1 _5051_ (.A1(_3303_),
    .A2(_3252_),
    .B1(_1455_),
    .C1(_1456_),
    .D1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__nand2_1 _5052_ (.A(_3273_),
    .B(_3177_),
    .Y(_1459_));
 sky130_fd_sc_hd__nand2_1 _5053_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1460_));
 sky130_fd_sc_hd__or2_1 _5054_ (.A(_0961_),
    .B(_3281_),
    .X(_1461_));
 sky130_fd_sc_hd__o2111a_1 _5055_ (.A1(_3183_),
    .A2(_3270_),
    .B1(_1459_),
    .C1(_1460_),
    .D1(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__or2_1 _5056_ (.A(_0658_),
    .B(_3294_),
    .X(_1463_));
 sky130_fd_sc_hd__o221a_1 _5057_ (.A1(_3279_),
    .A2(_3287_),
    .B1(_0653_),
    .B2(_3290_),
    .C1(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__o22ai_1 _5058_ (.A1(_0636_),
    .A2(_3305_),
    .B1(_0797_),
    .B2(_3308_),
    .Y(_1465_));
 sky130_fd_sc_hd__a221oi_1 _5059_ (.A1(_3214_),
    .A2(_3299_),
    .B1(_3205_),
    .B2(_3302_),
    .C1(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__and4_1 _5060_ (.A(_1458_),
    .B(_1462_),
    .C(_1464_),
    .D(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__inv_2 _5061_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1468_));
 sky130_fd_sc_hd__o22ai_1 _5062_ (.A1(_1346_),
    .A2(_3324_),
    .B1(_1468_),
    .B2(_3328_),
    .Y(_1469_));
 sky130_fd_sc_hd__a221oi_1 _5063_ (.A1(_3373_),
    .A2(_3317_),
    .B1(_0681_),
    .B2(_3321_),
    .C1(_1469_),
    .Y(_1470_));
 sky130_fd_sc_hd__nand2_1 _5064_ (.A(_3341_),
    .B(_0975_),
    .Y(_1471_));
 sky130_fd_sc_hd__nand2_1 _5065_ (.A(_3346_),
    .B(_0834_),
    .Y(_1472_));
 sky130_fd_sc_hd__nand2_1 _5066_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__a221oi_1 _5067_ (.A1(_1107_),
    .A2(_3334_),
    .B1(_3423_),
    .B2(_3338_),
    .C1(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _5068_ (.A(_3364_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1475_));
 sky130_fd_sc_hd__o21ai_1 _5069_ (.A1(_1097_),
    .A2(_3361_),
    .B1(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__a221oi_1 _5070_ (.A1(_3318_),
    .A2(_3354_),
    .B1(_3347_),
    .B2(_3358_),
    .C1(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1478_));
 sky130_fd_sc_hd__o21ai_1 _5072_ (.A1(_0686_),
    .A2(_3379_),
    .B1(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__a221oi_1 _5073_ (.A1(_3427_),
    .A2(_3372_),
    .B1(_3399_),
    .B2(_3376_),
    .C1(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__and4_1 _5074_ (.A(_1470_),
    .B(_1474_),
    .C(_1477_),
    .D(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__nand2_1 _5075_ (.A(_3393_),
    .B(_0322_),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2_1 _5076_ (.A(_3398_),
    .B(_0696_),
    .Y(_1483_));
 sky130_fd_sc_hd__or2_1 _5077_ (.A(_0985_),
    .B(_3403_),
    .X(_1484_));
 sky130_fd_sc_hd__o2111a_1 _5078_ (.A1(_0694_),
    .A2(_3390_),
    .B1(_1482_),
    .C1(_1483_),
    .D1(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__nand2_1 _5079_ (.A(_3411_),
    .B(_0853_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand2_1 _5080_ (.A(_3415_),
    .B(_0370_),
    .Y(_1487_));
 sky130_fd_sc_hd__or2_1 _5081_ (.A(_0364_),
    .B(_3420_),
    .X(_1488_));
 sky130_fd_sc_hd__o2111a_1 _5082_ (.A1(_0863_),
    .A2(_3408_),
    .B1(_1486_),
    .C1(_1487_),
    .D1(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_3436_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1490_));
 sky130_fd_sc_hd__o21ai_1 _5084_ (.A1(_3401_),
    .A2(_3433_),
    .B1(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__a221oi_1 _5085_ (.A1(_0980_),
    .A2(_3426_),
    .B1(_3416_),
    .B2(_3430_),
    .C1(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_0331_),
    .B(_0718_),
    .Y(_1493_));
 sky130_fd_sc_hd__o21ai_1 _5087_ (.A1(_0722_),
    .A2(_0328_),
    .B1(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__a221oi_1 _5088_ (.A1(_0360_),
    .A2(_3443_),
    .B1(_0380_),
    .B2(_0325_),
    .C1(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__and4_1 _5089_ (.A(_1485_),
    .B(_1489_),
    .C(_1492_),
    .D(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__and4_1 _5090_ (.A(_1454_),
    .B(_1467_),
    .C(_1481_),
    .D(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__inv_2 _5091_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1498_));
 sky130_fd_sc_hd__o22ai_1 _5092_ (.A1(_1376_),
    .A2(_0349_),
    .B1(_1498_),
    .B2(_0353_),
    .Y(_1499_));
 sky130_fd_sc_hd__a221oi_1 _5093_ (.A1(_0872_),
    .A2(_0342_),
    .B1(_0749_),
    .B2(_0346_),
    .C1(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_0369_),
    .B(_0868_),
    .Y(_1501_));
 sky130_fd_sc_hd__o21ai_1 _5095_ (.A1(_0374_),
    .A2(_0366_),
    .B1(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__a221oi_1 _5096_ (.A1(_0350_),
    .A2(_0359_),
    .B1(_0337_),
    .B2(_0363_),
    .C1(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__nand2_1 _5097_ (.A(_0379_),
    .B(_0343_),
    .Y(_1504_));
 sky130_fd_sc_hd__nand2_1 _5098_ (.A(_0384_),
    .B(_0403_),
    .Y(_1505_));
 sky130_fd_sc_hd__or2_1 _5099_ (.A(_0999_),
    .B(_0389_),
    .X(_1506_));
 sky130_fd_sc_hd__o2111a_1 _5100_ (.A1(_1253_),
    .A2(_0376_),
    .B1(_1504_),
    .C1(_1505_),
    .D1(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__nand2_1 _5101_ (.A(_0402_),
    .B(_0751_),
    .Y(_1508_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(_0407_),
    .B(_0500_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _5103_ (.A(_1508_),
    .B(_1509_),
    .Y(_1510_));
 sky130_fd_sc_hd__a221oi_1 _5104_ (.A1(_0897_),
    .A2(_0395_),
    .B1(_1032_),
    .B2(_0399_),
    .C1(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__and4_1 _5105_ (.A(_1500_),
    .B(_1503_),
    .C(_1507_),
    .D(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__o22ai_1 _5106_ (.A1(_0435_),
    .A2(_0423_),
    .B1(_0465_),
    .B2(_0426_),
    .Y(_1513_));
 sky130_fd_sc_hd__a221oi_1 _5107_ (.A1(_3122_),
    .A2(_0417_),
    .B1(_3125_),
    .B2(_0420_),
    .C1(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__nand2_1 _5108_ (.A(_0440_),
    .B(_0787_),
    .Y(_1515_));
 sky130_fd_sc_hd__o21ai_1 _5109_ (.A1(_3285_),
    .A2(_0437_),
    .B1(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__a221oi_1 _5110_ (.A1(_3129_),
    .A2(_0431_),
    .B1(_0625_),
    .B2(_0434_),
    .C1(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__nand2_1 _5111_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1518_));
 sky130_fd_sc_hd__o21ai_1 _5112_ (.A1(_0878_),
    .A2(_0452_),
    .B1(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__a221oi_1 _5113_ (.A1(_3110_),
    .A2(_0446_),
    .B1(_3113_),
    .B2(_0449_),
    .C1(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__o22ai_1 _5114_ (.A1(_3292_),
    .A2(_0467_),
    .B1(_0661_),
    .B2(_0470_),
    .Y(_1521_));
 sky130_fd_sc_hd__a221oi_2 _5115_ (.A1(_3246_),
    .A2(_0461_),
    .B1(_3256_),
    .B2(_0464_),
    .C1(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__and4_1 _5116_ (.A(_1514_),
    .B(_1517_),
    .C(_1520_),
    .D(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__o22ai_1 _5117_ (.A1(_0907_),
    .A2(_0487_),
    .B1(_1040_),
    .B2(_0490_),
    .Y(_1524_));
 sky130_fd_sc_hd__a221oi_1 _5118_ (.A1(_0569_),
    .A2(_0480_),
    .B1(_0580_),
    .B2(_0484_),
    .C1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nand2_1 _5119_ (.A(_0495_),
    .B(_0758_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_0499_),
    .B(_0474_),
    .Y(_1527_));
 sky130_fd_sc_hd__nand2_1 _5121_ (.A(_0504_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1528_));
 sky130_fd_sc_hd__nand2_1 _5122_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_1529_));
 sky130_fd_sc_hd__and4_1 _5123_ (.A(_1526_),
    .B(_1527_),
    .C(_1528_),
    .D(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__o22ai_1 _5124_ (.A1(_0893_),
    .A2(_0513_),
    .B1(_0533_),
    .B2(_0516_),
    .Y(_1531_));
 sky130_fd_sc_hd__a22o_1 _5125_ (.A1(_0519_),
    .A2(_0892_),
    .B1(_0521_),
    .B2(_0525_),
    .X(_1532_));
 sky130_fd_sc_hd__nor2_1 _5126_ (.A(_1531_),
    .B(_1532_),
    .Y(_1533_));
 sky130_fd_sc_hd__inv_2 _5127_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_1534_));
 sky130_fd_sc_hd__o22ai_1 _5128_ (.A1(_1412_),
    .A2(_0535_),
    .B1(_1534_),
    .B2(_0538_),
    .Y(_1535_));
 sky130_fd_sc_hd__a221oi_1 _5129_ (.A1(_0774_),
    .A2(_0528_),
    .B1(_0595_),
    .B2(_0532_),
    .C1(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__and4_1 _5130_ (.A(_1525_),
    .B(_1530_),
    .C(_1533_),
    .D(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__nand2_1 _5131_ (.A(_0555_),
    .B(_3072_),
    .Y(_1538_));
 sky130_fd_sc_hd__nand2_1 _5132_ (.A(_0560_),
    .B(_0924_),
    .Y(_1539_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(_1538_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__a221oi_1 _5134_ (.A1(_3084_),
    .A2(_0548_),
    .B1(_3087_),
    .B2(_0552_),
    .C1(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__nand2_1 _5135_ (.A(_0574_),
    .B(_0542_),
    .Y(_1542_));
 sky130_fd_sc_hd__nand2_1 _5136_ (.A(_0579_),
    .B(_0556_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _5137_ (.A(_1542_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__a221oi_1 _5138_ (.A1(_0776_),
    .A2(_0568_),
    .B1(_0561_),
    .B2(_0571_),
    .C1(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__inv_2 _5139_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1546_));
 sky130_fd_sc_hd__nand2_1 _5140_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1547_));
 sky130_fd_sc_hd__nand2_1 _5141_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1548_));
 sky130_fd_sc_hd__or2_1 _5142_ (.A(_1302_),
    .B(_0599_),
    .X(_1549_));
 sky130_fd_sc_hd__o2111a_1 _5143_ (.A1(_1546_),
    .A2(_0586_),
    .B1(_1547_),
    .C1(_1548_),
    .D1(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__nand2_1 _5144_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_1551_));
 sky130_fd_sc_hd__o21ai_1 _5145_ (.A1(_0731_),
    .A2(_0612_),
    .B1(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__a221oi_1 _5146_ (.A1(_3090_),
    .A2(_0605_),
    .B1(_3093_),
    .B2(_0609_),
    .C1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__and4_1 _5147_ (.A(_1541_),
    .B(_1545_),
    .C(_1550_),
    .D(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__and4_1 _5148_ (.A(_1512_),
    .B(_1523_),
    .C(_1537_),
    .D(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_0624_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_1556_));
 sky130_fd_sc_hd__nand3_1 _5150_ (.A(_1497_),
    .B(_1555_),
    .C(_1556_),
    .Y(_1557_));
 sky130_fd_sc_hd__nor2_1 _5151_ (.A(_3134_),
    .B(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__nor2_1 _5152_ (.A(_1437_),
    .B(_1558_),
    .Y(_0290_));
 sky130_fd_sc_hd__o21ai_1 _5153_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .A2(_3071_),
    .B1(_3132_),
    .Y(_1559_));
 sky130_fd_sc_hd__inv_2 _5154_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_3154_),
    .B(_3355_),
    .Y(_1561_));
 sky130_fd_sc_hd__a22o_1 _5156_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_1562_));
 sky130_fd_sc_hd__inv_2 _5157_ (.A(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__o211a_1 _5158_ (.A1(_1560_),
    .A2(_3147_),
    .B1(_1561_),
    .C1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_3190_),
    .B(_3167_),
    .Y(_1565_));
 sky130_fd_sc_hd__o21ai_1 _5160_ (.A1(_0792_),
    .A2(_3186_),
    .B1(_1565_),
    .Y(_1566_));
 sky130_fd_sc_hd__a221oi_1 _5161_ (.A1(_3135_),
    .A2(_3176_),
    .B1(_3155_),
    .B2(_3181_),
    .C1(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__nand2_1 _5162_ (.A(_3204_),
    .B(_3222_),
    .Y(_1568_));
 sky130_fd_sc_hd__nand2_1 _5163_ (.A(_3211_),
    .B(_3241_),
    .Y(_1569_));
 sky130_fd_sc_hd__or2_1 _5164_ (.A(_1193_),
    .B(_3219_),
    .X(_1570_));
 sky130_fd_sc_hd__o2111a_1 _5165_ (.A1(_1438_),
    .A2(_3200_),
    .B1(_1568_),
    .C1(_1569_),
    .D1(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__nand2_1 _5166_ (.A(_3234_),
    .B(_3325_),
    .Y(_1572_));
 sky130_fd_sc_hd__nand2_1 _5167_ (.A(_3240_),
    .B(_0677_),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2_1 _5168_ (.A(_1572_),
    .B(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__a221oi_1 _5169_ (.A1(_3312_),
    .A2(_3226_),
    .B1(_3318_),
    .B2(_3230_),
    .C1(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__and4_1 _5170_ (.A(_1564_),
    .B(_1567_),
    .C(_1571_),
    .D(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__nand2_1 _5171_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1577_));
 sky130_fd_sc_hd__nand2_1 _5172_ (.A(_3260_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1578_));
 sky130_fd_sc_hd__or2_1 _5173_ (.A(_0820_),
    .B(_3265_),
    .X(_1579_));
 sky130_fd_sc_hd__o2111a_1 _5174_ (.A1(_3306_),
    .A2(_3252_),
    .B1(_1577_),
    .C1(_1578_),
    .D1(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__nand2_1 _5175_ (.A(_3273_),
    .B(_3182_),
    .Y(_1581_));
 sky130_fd_sc_hd__nand2_1 _5176_ (.A(_3277_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1582_));
 sky130_fd_sc_hd__or2_1 _5177_ (.A(_1093_),
    .B(_3281_),
    .X(_1583_));
 sky130_fd_sc_hd__o2111a_1 _5178_ (.A1(_0636_),
    .A2(_3270_),
    .B1(_1581_),
    .C1(_1582_),
    .D1(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__or2_1 _5179_ (.A(_3268_),
    .B(_3294_),
    .X(_1585_));
 sky130_fd_sc_hd__o221a_1 _5180_ (.A1(_0658_),
    .A2(_3287_),
    .B1(_3279_),
    .B2(_3290_),
    .C1(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__o22ai_1 _5181_ (.A1(_0797_),
    .A2(_3305_),
    .B1(_3215_),
    .B2(_3308_),
    .Y(_1587_));
 sky130_fd_sc_hd__a221oi_1 _5182_ (.A1(_3205_),
    .A2(_3299_),
    .B1(_3195_),
    .B2(_3302_),
    .C1(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__and4_1 _5183_ (.A(_1580_),
    .B(_1584_),
    .C(_1586_),
    .D(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__inv_2 _5184_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1590_));
 sky130_fd_sc_hd__o22ai_1 _5185_ (.A1(_1468_),
    .A2(_3324_),
    .B1(_1590_),
    .B2(_3328_),
    .Y(_1591_));
 sky130_fd_sc_hd__a221oi_1 _5186_ (.A1(_0681_),
    .A2(_3317_),
    .B1(_0834_),
    .B2(_3321_),
    .C1(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__nand2_1 _5187_ (.A(_3341_),
    .B(_1107_),
    .Y(_1593_));
 sky130_fd_sc_hd__nand2_1 _5188_ (.A(_3346_),
    .B(_0975_),
    .Y(_1594_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(_1593_),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__a221oi_1 _5190_ (.A1(_3423_),
    .A2(_3334_),
    .B1(_3427_),
    .B2(_3338_),
    .C1(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _5191_ (.A(_3364_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_1597_));
 sky130_fd_sc_hd__o21ai_1 _5192_ (.A1(_1223_),
    .A2(_3361_),
    .B1(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__a221oi_1 _5193_ (.A1(_3347_),
    .A2(_3354_),
    .B1(_3342_),
    .B2(_3358_),
    .C1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__nand2_1 _5194_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1600_));
 sky130_fd_sc_hd__o21ai_1 _5195_ (.A1(_3401_),
    .A2(_3379_),
    .B1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__a221oi_1 _5196_ (.A1(_3399_),
    .A2(_3372_),
    .B1(_0689_),
    .B2(_3376_),
    .C1(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__and4_1 _5197_ (.A(_1592_),
    .B(_1596_),
    .C(_1599_),
    .D(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__nand2_1 _5198_ (.A(_3393_),
    .B(_0705_),
    .Y(_1604_));
 sky130_fd_sc_hd__nand2_1 _5199_ (.A(_3398_),
    .B(_3440_),
    .Y(_1605_));
 sky130_fd_sc_hd__or2_1 _5200_ (.A(_0326_),
    .B(_3403_),
    .X(_1606_));
 sky130_fd_sc_hd__o2111a_1 _5201_ (.A1(_0844_),
    .A2(_3390_),
    .B1(_1604_),
    .C1(_1605_),
    .D1(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__nand2_1 _5202_ (.A(_3411_),
    .B(_0854_),
    .Y(_1608_));
 sky130_fd_sc_hd__nand2_1 _5203_ (.A(_3415_),
    .B(_0356_),
    .Y(_1609_));
 sky130_fd_sc_hd__or2_1 _5204_ (.A(_0714_),
    .B(_3420_),
    .X(_1610_));
 sky130_fd_sc_hd__o2111a_1 _5205_ (.A1(_1002_),
    .A2(_3408_),
    .B1(_1608_),
    .C1(_1609_),
    .D1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_3436_),
    .B(_0980_),
    .Y(_1612_));
 sky130_fd_sc_hd__o21ai_1 _5207_ (.A1(_0691_),
    .A2(_3433_),
    .B1(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__a221oi_1 _5208_ (.A1(_3416_),
    .A2(_3426_),
    .B1(_0696_),
    .B2(_3430_),
    .C1(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__nand2_1 _5209_ (.A(_0331_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1615_));
 sky130_fd_sc_hd__o21ai_1 _5210_ (.A1(_0374_),
    .A2(_0328_),
    .B1(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__a221oi_1 _5211_ (.A1(_0380_),
    .A2(_3443_),
    .B1(_0718_),
    .B2(_0325_),
    .C1(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__and4_1 _5212_ (.A(_1607_),
    .B(_1611_),
    .C(_1614_),
    .D(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__and4_1 _5213_ (.A(_1576_),
    .B(_1589_),
    .C(_1603_),
    .D(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__inv_2 _5214_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1620_));
 sky130_fd_sc_hd__o22ai_1 _5215_ (.A1(_1498_),
    .A2(_0349_),
    .B1(_1620_),
    .B2(_0353_),
    .Y(_1621_));
 sky130_fd_sc_hd__a221oi_1 _5216_ (.A1(_0749_),
    .A2(_0342_),
    .B1(_0500_),
    .B2(_0346_),
    .C1(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__nand2_1 _5217_ (.A(_0369_),
    .B(_0350_),
    .Y(_1623_));
 sky130_fd_sc_hd__o21ai_1 _5218_ (.A1(_0347_),
    .A2(_0366_),
    .B1(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__a221oi_1 _5219_ (.A1(_0337_),
    .A2(_0359_),
    .B1(_0343_),
    .B2(_0363_),
    .C1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(_0379_),
    .B(_0408_),
    .Y(_1626_));
 sky130_fd_sc_hd__nand2_1 _5221_ (.A(_0384_),
    .B(_0392_),
    .Y(_1627_));
 sky130_fd_sc_hd__or2_1 _5222_ (.A(_1129_),
    .B(_0389_),
    .X(_1628_));
 sky130_fd_sc_hd__o2111a_1 _5223_ (.A1(_1376_),
    .A2(_0376_),
    .B1(_1626_),
    .C1(_1627_),
    .D1(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__nand2_1 _5224_ (.A(_0402_),
    .B(_0897_),
    .Y(_1630_));
 sky130_fd_sc_hd__nand2_1 _5225_ (.A(_0407_),
    .B(_0751_),
    .Y(_1631_));
 sky130_fd_sc_hd__nand2_1 _5226_ (.A(_1630_),
    .B(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__a221oi_1 _5227_ (.A1(_1032_),
    .A2(_0395_),
    .B1(_0522_),
    .B2(_0399_),
    .C1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__and4_1 _5228_ (.A(_1622_),
    .B(_1625_),
    .C(_1629_),
    .D(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__o22ai_1 _5229_ (.A1(_0465_),
    .A2(_0423_),
    .B1(_0468_),
    .B2(_0426_),
    .Y(_1635_));
 sky130_fd_sc_hd__a221oi_1 _5230_ (.A1(_3125_),
    .A2(_0417_),
    .B1(_3129_),
    .B2(_0420_),
    .C1(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _5231_ (.A(_0440_),
    .B(_3284_),
    .Y(_1637_));
 sky130_fd_sc_hd__o21ai_1 _5232_ (.A1(_3292_),
    .A2(_0437_),
    .B1(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__a221oi_1 _5233_ (.A1(_0625_),
    .A2(_0431_),
    .B1(_0787_),
    .B2(_0434_),
    .C1(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1640_));
 sky130_fd_sc_hd__o21ai_1 _5235_ (.A1(_1015_),
    .A2(_0452_),
    .B1(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__a221oi_1 _5236_ (.A1(_3113_),
    .A2(_0446_),
    .B1(_3116_),
    .B2(_0449_),
    .C1(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__o22ai_1 _5237_ (.A1(_0661_),
    .A2(_0467_),
    .B1(_3247_),
    .B2(_0470_),
    .Y(_1643_));
 sky130_fd_sc_hd__a221oi_1 _5238_ (.A1(_3256_),
    .A2(_0461_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .B2(_0464_),
    .C1(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__and4_1 _5239_ (.A(_1636_),
    .B(_1639_),
    .C(_1642_),
    .D(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__o22ai_1 _5240_ (.A1(_1040_),
    .A2(_0487_),
    .B1(_1167_),
    .B2(_0490_),
    .Y(_1646_));
 sky130_fd_sc_hd__a221oi_1 _5241_ (.A1(_0580_),
    .A2(_0480_),
    .B1(_0575_),
    .B2(_0484_),
    .C1(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_0495_),
    .B(_0904_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_0499_),
    .B(_0481_),
    .Y(_1649_));
 sky130_fd_sc_hd__nand2_1 _5244_ (.A(_0504_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1650_));
 sky130_fd_sc_hd__nand2_1 _5245_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_1651_));
 sky130_fd_sc_hd__and4_1 _5246_ (.A(_1648_),
    .B(_1649_),
    .C(_1650_),
    .D(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__o22ai_1 _5247_ (.A1(_0533_),
    .A2(_0513_),
    .B1(_0536_),
    .B2(_0516_),
    .Y(_1653_));
 sky130_fd_sc_hd__a22o_1 _5248_ (.A1(_0519_),
    .A2(_0525_),
    .B1(_0521_),
    .B2(_0529_),
    .X(_1654_));
 sky130_fd_sc_hd__nor2_1 _5249_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__o22ai_1 _5250_ (.A1(_1534_),
    .A2(_0535_),
    .B1(_0597_),
    .B2(_0538_),
    .Y(_1656_));
 sky130_fd_sc_hd__a221oi_1 _5251_ (.A1(_0595_),
    .A2(_0528_),
    .B1(_0776_),
    .B2(_0532_),
    .C1(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__and4_1 _5252_ (.A(_1647_),
    .B(_1652_),
    .C(_1655_),
    .D(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__nand2_1 _5253_ (.A(_0555_),
    .B(_3084_),
    .Y(_1659_));
 sky130_fd_sc_hd__nand2_1 _5254_ (.A(_0560_),
    .B(_3072_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand2_1 _5255_ (.A(_1659_),
    .B(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__a221oi_1 _5256_ (.A1(_3087_),
    .A2(_0548_),
    .B1(_3090_),
    .B2(_0552_),
    .C1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__nand2_1 _5257_ (.A(_0574_),
    .B(_0549_),
    .Y(_1663_));
 sky130_fd_sc_hd__nand2_1 _5258_ (.A(_0579_),
    .B(_0542_),
    .Y(_1664_));
 sky130_fd_sc_hd__nand2_1 _5259_ (.A(_1663_),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__a221oi_1 _5260_ (.A1(_0561_),
    .A2(_0568_),
    .B1(_0556_),
    .B2(_0571_),
    .C1(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__nand2_1 _5261_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1667_));
 sky130_fd_sc_hd__nand2_1 _5262_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1668_));
 sky130_fd_sc_hd__or2_1 _5263_ (.A(_1424_),
    .B(_0599_),
    .X(_1669_));
 sky130_fd_sc_hd__o2111a_1 _5264_ (.A1(_0610_),
    .A2(_0586_),
    .B1(_1667_),
    .C1(_1668_),
    .D1(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1671_));
 sky130_fd_sc_hd__o21ai_1 _5266_ (.A1(_0878_),
    .A2(_0612_),
    .B1(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__a221oi_1 _5267_ (.A1(_3093_),
    .A2(_0605_),
    .B1(_3098_),
    .B2(_0609_),
    .C1(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__and4_1 _5268_ (.A(_1662_),
    .B(_1666_),
    .C(_1670_),
    .D(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__and4_1 _5269_ (.A(_1634_),
    .B(_1645_),
    .C(_1658_),
    .D(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__nand2_1 _5270_ (.A(_0624_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_1676_));
 sky130_fd_sc_hd__nand3_1 _5271_ (.A(_1619_),
    .B(_1675_),
    .C(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__nor2_1 _5272_ (.A(_3134_),
    .B(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__nor2_1 _5273_ (.A(_1559_),
    .B(_1678_),
    .Y(_0289_));
 sky130_fd_sc_hd__o21ai_1 _5274_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .A2(_3070_),
    .B1(_3132_),
    .Y(_1679_));
 sky130_fd_sc_hd__inv_2 _5275_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_1680_));
 sky130_fd_sc_hd__nand2_1 _5276_ (.A(_3154_),
    .B(_0675_),
    .Y(_1681_));
 sky130_fd_sc_hd__a22o_1 _5277_ (.A1(_3161_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .B1(_3166_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_1682_));
 sky130_fd_sc_hd__inv_2 _5278_ (.A(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__o211a_1 _5279_ (.A1(_1680_),
    .A2(_3147_),
    .B1(_1681_),
    .C1(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__nand2_1 _5280_ (.A(_3190_),
    .B(_3241_),
    .Y(_1685_));
 sky130_fd_sc_hd__o21ai_1 _5281_ (.A1(_0934_),
    .A2(_3186_),
    .B1(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__a221oi_1 _5282_ (.A1(_3155_),
    .A2(_3176_),
    .B1(_0631_),
    .B2(_3181_),
    .C1(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__nand2_1 _5283_ (.A(_3204_),
    .B(_3227_),
    .Y(_1688_));
 sky130_fd_sc_hd__nand2_1 _5284_ (.A(_3211_),
    .B(_3235_),
    .Y(_1689_));
 sky130_fd_sc_hd__or2_1 _5285_ (.A(_1316_),
    .B(_3219_),
    .X(_1690_));
 sky130_fd_sc_hd__o2111a_1 _5286_ (.A1(_1560_),
    .A2(_3200_),
    .B1(_1688_),
    .C1(_1689_),
    .D1(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__nand2_1 _5287_ (.A(_3234_),
    .B(_3312_),
    .Y(_1692_));
 sky130_fd_sc_hd__nand2_1 _5288_ (.A(_3240_),
    .B(_3325_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_1 _5289_ (.A(_1692_),
    .B(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__a221oi_1 _5290_ (.A1(_3318_),
    .A2(_3226_),
    .B1(_3347_),
    .B2(_3230_),
    .C1(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__and4_1 _5291_ (.A(_1684_),
    .B(_1687_),
    .C(_1691_),
    .D(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__nand2_1 _5292_ (.A(_3255_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1697_));
 sky130_fd_sc_hd__nand2_1 _5293_ (.A(_3260_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_1698_));
 sky130_fd_sc_hd__or2_1 _5294_ (.A(_0961_),
    .B(_3265_),
    .X(_1699_));
 sky130_fd_sc_hd__o2111a_1 _5295_ (.A1(_0664_),
    .A2(_3252_),
    .B1(_1697_),
    .C1(_1698_),
    .D1(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__nand2_1 _5296_ (.A(_3273_),
    .B(_3191_),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _5297_ (.A(_3277_),
    .B(_3177_),
    .Y(_1702_));
 sky130_fd_sc_hd__or2_1 _5298_ (.A(_3183_),
    .B(_3281_),
    .X(_1703_));
 sky130_fd_sc_hd__o2111a_1 _5299_ (.A1(_0797_),
    .A2(_3270_),
    .B1(_1701_),
    .C1(_1702_),
    .D1(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__or2_1 _5300_ (.A(_3303_),
    .B(_3294_),
    .X(_1705_));
 sky130_fd_sc_hd__o221a_1 _5301_ (.A1(_3268_),
    .A2(_3287_),
    .B1(_0658_),
    .B2(_3290_),
    .C1(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__o22ai_1 _5302_ (.A1(_3215_),
    .A2(_3305_),
    .B1(_0642_),
    .B2(_3308_),
    .Y(_1707_));
 sky130_fd_sc_hd__a221oi_1 _5303_ (.A1(_3195_),
    .A2(_3299_),
    .B1(_3135_),
    .B2(_3302_),
    .C1(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__and4_1 _5304_ (.A(_1700_),
    .B(_1704_),
    .C(_1706_),
    .D(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__inv_2 _5305_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1710_));
 sky130_fd_sc_hd__o22ai_1 _5306_ (.A1(_1590_),
    .A2(_3324_),
    .B1(_1710_),
    .B2(_3328_),
    .Y(_1711_));
 sky130_fd_sc_hd__a221oi_1 _5307_ (.A1(_0834_),
    .A2(_3317_),
    .B1(_0975_),
    .B2(_3321_),
    .C1(_1711_),
    .Y(_1712_));
 sky130_fd_sc_hd__nand2_1 _5308_ (.A(_3341_),
    .B(_3423_),
    .Y(_1713_));
 sky130_fd_sc_hd__nand2_1 _5309_ (.A(_3346_),
    .B(_1107_),
    .Y(_1714_));
 sky130_fd_sc_hd__nand2_1 _5310_ (.A(_1713_),
    .B(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__a221oi_1 _5311_ (.A1(_3427_),
    .A2(_3334_),
    .B1(_3399_),
    .B2(_3338_),
    .C1(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__nand2_1 _5312_ (.A(_3364_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1717_));
 sky130_fd_sc_hd__o21ai_1 _5313_ (.A1(_1346_),
    .A2(_3361_),
    .B1(_1717_),
    .Y(_1718_));
 sky130_fd_sc_hd__a221oi_1 _5314_ (.A1(_3342_),
    .A2(_3354_),
    .B1(_3331_),
    .B2(_3358_),
    .C1(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__nand2_1 _5315_ (.A(_3382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1720_));
 sky130_fd_sc_hd__o21ai_1 _5316_ (.A1(_0691_),
    .A2(_3379_),
    .B1(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__a221oi_1 _5317_ (.A1(_0689_),
    .A2(_3372_),
    .B1(_3394_),
    .B2(_3376_),
    .C1(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__and4_1 _5318_ (.A(_1712_),
    .B(_1716_),
    .C(_1719_),
    .D(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__nand2_1 _5319_ (.A(_3393_),
    .B(_0853_),
    .Y(_1724_));
 sky130_fd_sc_hd__nand2_1 _5320_ (.A(_3398_),
    .B(_0322_),
    .Y(_1725_));
 sky130_fd_sc_hd__or2_1 _5321_ (.A(_0364_),
    .B(_3403_),
    .X(_1726_));
 sky130_fd_sc_hd__o2111a_1 _5322_ (.A1(_0985_),
    .A2(_3390_),
    .B1(_1724_),
    .C1(_1725_),
    .D1(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__nand2_1 _5323_ (.A(_3411_),
    .B(_0370_),
    .Y(_1728_));
 sky130_fd_sc_hd__nand2_1 _5324_ (.A(_3415_),
    .B(_0360_),
    .Y(_1729_));
 sky130_fd_sc_hd__or2_1 _5325_ (.A(_0863_),
    .B(_3420_),
    .X(_1730_));
 sky130_fd_sc_hd__o2111a_1 _5326_ (.A1(_1132_),
    .A2(_3408_),
    .B1(_1728_),
    .C1(_1729_),
    .D1(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__nand2_1 _5327_ (.A(_3436_),
    .B(_3416_),
    .Y(_1732_));
 sky130_fd_sc_hd__o21ai_1 _5328_ (.A1(_3418_),
    .A2(_3433_),
    .B1(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__a221oi_1 _5329_ (.A1(_0696_),
    .A2(_3426_),
    .B1(_3440_),
    .B2(_3430_),
    .C1(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _5330_ (.A(_0331_),
    .B(_0720_),
    .Y(_1735_));
 sky130_fd_sc_hd__o21ai_1 _5331_ (.A1(_0347_),
    .A2(_0328_),
    .B1(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__a221oi_1 _5332_ (.A1(_0718_),
    .A2(_3443_),
    .B1(_0385_),
    .B2(_0325_),
    .C1(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__and4_1 _5333_ (.A(_1727_),
    .B(_1731_),
    .C(_1734_),
    .D(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__and4_1 _5334_ (.A(_1696_),
    .B(_1709_),
    .C(_1723_),
    .D(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__inv_2 _5335_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1740_));
 sky130_fd_sc_hd__o22ai_1 _5336_ (.A1(_1620_),
    .A2(_0349_),
    .B1(_1740_),
    .B2(_0353_),
    .Y(_1741_));
 sky130_fd_sc_hd__a221oi_1 _5337_ (.A1(_0500_),
    .A2(_0342_),
    .B1(_0751_),
    .B2(_0346_),
    .C1(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__nand2_1 _5338_ (.A(_0369_),
    .B(_0337_),
    .Y(_1743_));
 sky130_fd_sc_hd__o21ai_1 _5339_ (.A1(_0351_),
    .A2(_0366_),
    .B1(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__a221oi_1 _5340_ (.A1(_0343_),
    .A2(_0359_),
    .B1(_0408_),
    .B2(_0363_),
    .C1(_1744_),
    .Y(_1745_));
 sky130_fd_sc_hd__nand2_1 _5341_ (.A(_0379_),
    .B(_0403_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5342_ (.A(_0384_),
    .B(_0396_),
    .Y(_1747_));
 sky130_fd_sc_hd__or2_1 _5343_ (.A(_1253_),
    .B(_0389_),
    .X(_1748_));
 sky130_fd_sc_hd__o2111a_1 _5344_ (.A1(_1498_),
    .A2(_0376_),
    .B1(_1746_),
    .C1(_1747_),
    .D1(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__nand2_1 _5345_ (.A(_0402_),
    .B(_1032_),
    .Y(_1750_));
 sky130_fd_sc_hd__nand2_1 _5346_ (.A(_0407_),
    .B(_0897_),
    .Y(_1751_));
 sky130_fd_sc_hd__nand2_1 _5347_ (.A(_1750_),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__a221oi_1 _5348_ (.A1(_0522_),
    .A2(_0395_),
    .B1(_0758_),
    .B2(_0399_),
    .C1(_1752_),
    .Y(_1753_));
 sky130_fd_sc_hd__and4_1 _5349_ (.A(_1742_),
    .B(_1745_),
    .C(_1749_),
    .D(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__o22ai_1 _5350_ (.A1(_0468_),
    .A2(_0423_),
    .B1(_0741_),
    .B2(_0426_),
    .Y(_1755_));
 sky130_fd_sc_hd__a221oi_1 _5351_ (.A1(_3129_),
    .A2(_0417_),
    .B1(_0625_),
    .B2(_0420_),
    .C1(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _5352_ (.A(_0440_),
    .B(_3291_),
    .Y(_1757_));
 sky130_fd_sc_hd__o21ai_1 _5353_ (.A1(_0661_),
    .A2(_0437_),
    .B1(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__a221oi_1 _5354_ (.A1(_0787_),
    .A2(_0431_),
    .B1(_3284_),
    .B2(_0434_),
    .C1(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1760_));
 sky130_fd_sc_hd__o21ai_1 _5356_ (.A1(_1145_),
    .A2(_0452_),
    .B1(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__a221oi_1 _5357_ (.A1(_3116_),
    .A2(_0446_),
    .B1(_3119_),
    .B2(_0449_),
    .C1(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__o22ai_1 _5358_ (.A1(_3247_),
    .A2(_0467_),
    .B1(_0650_),
    .B2(_0470_),
    .Y(_1763_));
 sky130_fd_sc_hd__a221oi_1 _5359_ (.A1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .A2(_0461_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .B2(_0464_),
    .C1(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__and4_1 _5360_ (.A(_1756_),
    .B(_1759_),
    .C(_1762_),
    .D(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__o22ai_1 _5361_ (.A1(_1167_),
    .A2(_0487_),
    .B1(_1290_),
    .B2(_0490_),
    .Y(_1766_));
 sky130_fd_sc_hd__a221oi_1 _5362_ (.A1(_0575_),
    .A2(_0480_),
    .B1(_0590_),
    .B2(_0484_),
    .C1(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__nand2_1 _5363_ (.A(_0495_),
    .B(_0474_),
    .Y(_1768_));
 sky130_fd_sc_hd__nand2_1 _5364_ (.A(_0499_),
    .B(_0745_),
    .Y(_1769_));
 sky130_fd_sc_hd__nand2_1 _5365_ (.A(_0504_),
    .B(_0904_),
    .Y(_1770_));
 sky130_fd_sc_hd__nand2_1 _5366_ (.A(_0508_),
    .B(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_1771_));
 sky130_fd_sc_hd__and4_1 _5367_ (.A(_1768_),
    .B(_1769_),
    .C(_1770_),
    .D(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__o22ai_1 _5368_ (.A1(_0536_),
    .A2(_0513_),
    .B1(_0761_),
    .B2(_0516_),
    .Y(_1773_));
 sky130_fd_sc_hd__a22o_1 _5369_ (.A1(_0519_),
    .A2(_0529_),
    .B1(_0521_),
    .B2(_0565_),
    .X(_1774_));
 sky130_fd_sc_hd__nor2_1 _5370_ (.A(_1773_),
    .B(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__o22ai_1 _5371_ (.A1(_0597_),
    .A2(_0535_),
    .B1(_0778_),
    .B2(_0538_),
    .Y(_1776_));
 sky130_fd_sc_hd__a221oi_1 _5372_ (.A1(_0776_),
    .A2(_0528_),
    .B1(_0561_),
    .B2(_0532_),
    .C1(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__and4_1 _5373_ (.A(_1767_),
    .B(_1772_),
    .C(_1775_),
    .D(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__nand2_1 _5374_ (.A(_0555_),
    .B(_3087_),
    .Y(_1779_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(_0560_),
    .B(_3084_),
    .Y(_1780_));
 sky130_fd_sc_hd__nand2_1 _5376_ (.A(_1779_),
    .B(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__a221oi_1 _5377_ (.A1(_3090_),
    .A2(_0548_),
    .B1(_3093_),
    .B2(_0552_),
    .C1(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(_0574_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1783_));
 sky130_fd_sc_hd__nand2_1 _5379_ (.A(_0579_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1784_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(_1783_),
    .B(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__a221oi_1 _5381_ (.A1(_0556_),
    .A2(_0568_),
    .B1(_0542_),
    .B2(_0571_),
    .C1(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__nand2_1 _5382_ (.A(_0589_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1787_));
 sky130_fd_sc_hd__nand2_1 _5383_ (.A(_0594_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_1788_));
 sky130_fd_sc_hd__or2_1 _5384_ (.A(_1546_),
    .B(_0599_),
    .X(_1789_));
 sky130_fd_sc_hd__o2111a_1 _5385_ (.A1(_0450_),
    .A2(_0586_),
    .B1(_1787_),
    .C1(_1788_),
    .D1(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__nand2_1 _5386_ (.A(_0615_),
    .B(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_1791_));
 sky130_fd_sc_hd__o21ai_1 _5387_ (.A1(_1015_),
    .A2(_0612_),
    .B1(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__a221oi_1 _5388_ (.A1(_3098_),
    .A2(_0605_),
    .B1(_3101_),
    .B2(_0609_),
    .C1(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__and4_1 _5389_ (.A(_1782_),
    .B(_1786_),
    .C(_1790_),
    .D(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__and4_1 _5390_ (.A(_1754_),
    .B(_1765_),
    .C(_1778_),
    .D(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__nand2_1 _5391_ (.A(_0624_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_1796_));
 sky130_fd_sc_hd__nand3_1 _5392_ (.A(_1739_),
    .B(_1795_),
    .C(_1796_),
    .Y(_1797_));
 sky130_fd_sc_hd__nor2_1 _5393_ (.A(_3134_),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__nor2_1 _5394_ (.A(_1679_),
    .B(_1798_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21ai_1 _5395_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .A2(_3070_),
    .B1(_3009_),
    .Y(_1799_));
 sky130_fd_sc_hd__nand2_1 _5396_ (.A(_3153_),
    .B(_3365_),
    .Y(_1800_));
 sky130_fd_sc_hd__a22o_1 _5397_ (.A1(_3160_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .B1(_3165_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_1801_));
 sky130_fd_sc_hd__inv_2 _5398_ (.A(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__o211a_1 _5399_ (.A1(_3359_),
    .A2(_3146_),
    .B1(_1800_),
    .C1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__nand2_1 _5400_ (.A(_3189_),
    .B(_3235_),
    .Y(_1804_));
 sky130_fd_sc_hd__o21ai_1 _5401_ (.A1(_1066_),
    .A2(_3185_),
    .B1(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__a221oi_1 _5402_ (.A1(_0631_),
    .A2(_3175_),
    .B1(_3167_),
    .B2(_3180_),
    .C1(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _5403_ (.A(_3203_),
    .B(_3351_),
    .Y(_1807_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(_3210_),
    .B(_3222_),
    .Y(_1808_));
 sky130_fd_sc_hd__or2_1 _5405_ (.A(_1438_),
    .B(_3218_),
    .X(_1809_));
 sky130_fd_sc_hd__o2111a_1 _5406_ (.A1(_1680_),
    .A2(_3199_),
    .B1(_1807_),
    .C1(_1808_),
    .D1(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__nand2_1 _5407_ (.A(_3233_),
    .B(_3318_),
    .Y(_1811_));
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_3239_),
    .B(_3312_),
    .Y(_1812_));
 sky130_fd_sc_hd__nand2_1 _5409_ (.A(_1811_),
    .B(_1812_),
    .Y(_1813_));
 sky130_fd_sc_hd__a221oi_1 _5410_ (.A1(_3347_),
    .A2(_3225_),
    .B1(_3342_),
    .B2(_3229_),
    .C1(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__and4_1 _5411_ (.A(_1803_),
    .B(_1806_),
    .C(_1810_),
    .D(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__nand2_1 _5412_ (.A(_3254_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1816_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(_3259_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_1817_));
 sky130_fd_sc_hd__or2_1 _5414_ (.A(_1093_),
    .B(_3264_),
    .X(_1818_));
 sky130_fd_sc_hd__o2111a_1 _5415_ (.A1(_0820_),
    .A2(_3251_),
    .B1(_1816_),
    .C1(_1817_),
    .D1(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__nand2_1 _5416_ (.A(_3272_),
    .B(_3212_),
    .Y(_1820_));
 sky130_fd_sc_hd__nand2_1 _5417_ (.A(_3276_),
    .B(_3182_),
    .Y(_1821_));
 sky130_fd_sc_hd__or2_1 _5418_ (.A(_0636_),
    .B(_3280_),
    .X(_1822_));
 sky130_fd_sc_hd__o2111a_1 _5419_ (.A1(_3215_),
    .A2(_3269_),
    .B1(_1820_),
    .C1(_1821_),
    .D1(_1822_),
    .X(_1823_));
 sky130_fd_sc_hd__or2_1 _5420_ (.A(_3306_),
    .B(_3293_),
    .X(_1824_));
 sky130_fd_sc_hd__o221a_1 _5421_ (.A1(_3303_),
    .A2(_3286_),
    .B1(_3268_),
    .B2(_3289_),
    .C1(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__o22ai_1 _5422_ (.A1(_0642_),
    .A2(_3304_),
    .B1(_3196_),
    .B2(_3307_),
    .Y(_1826_));
 sky130_fd_sc_hd__a221oi_1 _5423_ (.A1(_3135_),
    .A2(_3298_),
    .B1(_3155_),
    .B2(_3301_),
    .C1(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__and4_1 _5424_ (.A(_1819_),
    .B(_1823_),
    .C(_1825_),
    .D(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__o22ai_1 _5425_ (.A1(_1710_),
    .A2(_3323_),
    .B1(_3377_),
    .B2(_3327_),
    .Y(_1829_));
 sky130_fd_sc_hd__a221oi_1 _5426_ (.A1(_0975_),
    .A2(_3316_),
    .B1(_1107_),
    .B2(_3320_),
    .C1(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_3340_),
    .B(_3427_),
    .Y(_1831_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_3345_),
    .B(_3423_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1831_),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__a221oi_1 _5430_ (.A1(_3399_),
    .A2(_3333_),
    .B1(_0689_),
    .B2(_3337_),
    .C1(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_3363_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1835_));
 sky130_fd_sc_hd__o21ai_1 _5432_ (.A1(_1468_),
    .A2(_3360_),
    .B1(_1835_),
    .Y(_1836_));
 sky130_fd_sc_hd__a221oi_1 _5433_ (.A1(_3331_),
    .A2(_3353_),
    .B1(_3335_),
    .B2(_3357_),
    .C1(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__nand2_1 _5434_ (.A(_3381_),
    .B(_0839_),
    .Y(_1838_));
 sky130_fd_sc_hd__o21ai_1 _5435_ (.A1(_3418_),
    .A2(_3378_),
    .B1(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__a221oi_1 _5436_ (.A1(_3394_),
    .A2(_3371_),
    .B1(_0687_),
    .B2(_3375_),
    .C1(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__and4_1 _5437_ (.A(_1830_),
    .B(_1834_),
    .C(_1837_),
    .D(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(_3392_),
    .B(_0854_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _5439_ (.A(_3397_),
    .B(_0705_),
    .Y(_1843_));
 sky130_fd_sc_hd__or2_1 _5440_ (.A(_0714_),
    .B(_3402_),
    .X(_1844_));
 sky130_fd_sc_hd__o2111a_1 _5441_ (.A1(_0326_),
    .A2(_3389_),
    .B1(_1842_),
    .C1(_1843_),
    .D1(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_3410_),
    .B(_0356_),
    .Y(_1846_));
 sky130_fd_sc_hd__nand2_1 _5443_ (.A(_3414_),
    .B(_0380_),
    .Y(_1847_));
 sky130_fd_sc_hd__or2_1 _5444_ (.A(_1002_),
    .B(_3419_),
    .X(_1848_));
 sky130_fd_sc_hd__o2111a_1 _5445_ (.A1(_0387_),
    .A2(_3407_),
    .B1(_1846_),
    .C1(_1847_),
    .D1(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__nand2_1 _5446_ (.A(_3435_),
    .B(_0696_),
    .Y(_1850_));
 sky130_fd_sc_hd__o21ai_1 _5447_ (.A1(_0698_),
    .A2(_3432_),
    .B1(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__a221oi_1 _5448_ (.A1(_3440_),
    .A2(_3425_),
    .B1(_0322_),
    .B2(_3429_),
    .C1(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__nand2_1 _5449_ (.A(_0330_),
    .B(_0868_),
    .Y(_1853_));
 sky130_fd_sc_hd__o21ai_1 _5450_ (.A1(_0351_),
    .A2(_0327_),
    .B1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__a221oi_1 _5451_ (.A1(_0385_),
    .A2(_3442_),
    .B1(_0720_),
    .B2(_0324_),
    .C1(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__and4_1 _5452_ (.A(_1845_),
    .B(_1849_),
    .C(_1852_),
    .D(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__and4_1 _5453_ (.A(_1815_),
    .B(_1828_),
    .C(_1841_),
    .D(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__inv_2 _5454_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1858_));
 sky130_fd_sc_hd__o22ai_1 _5455_ (.A1(_1740_),
    .A2(_0348_),
    .B1(_1858_),
    .B2(_0352_),
    .Y(_1859_));
 sky130_fd_sc_hd__a221oi_1 _5456_ (.A1(_0751_),
    .A2(_0341_),
    .B1(_0897_),
    .B2(_0345_),
    .C1(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(_0368_),
    .B(_0343_),
    .Y(_1861_));
 sky130_fd_sc_hd__o21ai_1 _5458_ (.A1(_0711_),
    .A2(_0365_),
    .B1(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__a221oi_1 _5459_ (.A1(_0408_),
    .A2(_0358_),
    .B1(_0403_),
    .B2(_0362_),
    .C1(_1862_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand2_1 _5460_ (.A(_0378_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1864_));
 sky130_fd_sc_hd__nand2_1 _5461_ (.A(_0383_),
    .B(_0725_),
    .Y(_1865_));
 sky130_fd_sc_hd__or2_1 _5462_ (.A(_1376_),
    .B(_0388_),
    .X(_1866_));
 sky130_fd_sc_hd__o2111a_1 _5463_ (.A1(_1620_),
    .A2(_0375_),
    .B1(_1864_),
    .C1(_1865_),
    .D1(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__nand2_1 _5464_ (.A(_0401_),
    .B(_0522_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_0406_),
    .B(_1032_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _5466_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__a221oi_1 _5467_ (.A1(_0758_),
    .A2(_0394_),
    .B1(_0904_),
    .B2(_0398_),
    .C1(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__and4_1 _5468_ (.A(_1860_),
    .B(_1863_),
    .C(_1867_),
    .D(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__o22ai_1 _5469_ (.A1(_0741_),
    .A2(_0422_),
    .B1(_0888_),
    .B2(_0425_),
    .Y(_1873_));
 sky130_fd_sc_hd__a221oi_1 _5470_ (.A1(_0625_),
    .A2(_0416_),
    .B1(_0787_),
    .B2(_0419_),
    .C1(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__nand2_1 _5471_ (.A(_0439_),
    .B(_3261_),
    .Y(_1875_));
 sky130_fd_sc_hd__o21ai_1 _5472_ (.A1(_3247_),
    .A2(_0436_),
    .B1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__a221oi_1 _5473_ (.A1(_3284_),
    .A2(_0430_),
    .B1(_3291_),
    .B2(_0433_),
    .C1(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _5474_ (.A(_0454_),
    .B(_3116_),
    .Y(_1878_));
 sky130_fd_sc_hd__o21ai_1 _5475_ (.A1(_1268_),
    .A2(_0451_),
    .B1(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hd__a221oi_1 _5476_ (.A1(_3119_),
    .A2(_0445_),
    .B1(_3122_),
    .B2(_0448_),
    .C1(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__o22ai_1 _5477_ (.A1(_0650_),
    .A2(_0466_),
    .B1(_3263_),
    .B2(_0469_),
    .Y(_1881_));
 sky130_fd_sc_hd__a221oi_1 _5478_ (.A1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .A2(_0460_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .B2(_0463_),
    .C1(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__and4_1 _5479_ (.A(_1874_),
    .B(_1877_),
    .C(_1880_),
    .D(_1882_),
    .X(_1883_));
 sky130_fd_sc_hd__o22ai_1 _5480_ (.A1(_1290_),
    .A2(_0486_),
    .B1(_1412_),
    .B2(_0489_),
    .Y(_1884_));
 sky130_fd_sc_hd__a221oi_1 _5481_ (.A1(_0590_),
    .A2(_0479_),
    .B1(_0774_),
    .B2(_0483_),
    .C1(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_0494_),
    .B(_0481_),
    .Y(_1886_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_0498_),
    .B(_0892_),
    .Y(_1887_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_0503_),
    .B(_0474_),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_1 _5485_ (.A(_0507_),
    .B(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_1889_));
 sky130_fd_sc_hd__and4_1 _5486_ (.A(_1886_),
    .B(_1887_),
    .C(_1888_),
    .D(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__o22ai_1 _5487_ (.A1(_0761_),
    .A2(_0512_),
    .B1(_0907_),
    .B2(_0515_),
    .Y(_1891_));
 sky130_fd_sc_hd__a22o_1 _5488_ (.A1(_0518_),
    .A2(_0565_),
    .B1(_0520_),
    .B2(_0569_),
    .X(_1892_));
 sky130_fd_sc_hd__nor2_1 _5489_ (.A(_1891_),
    .B(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__o22ai_1 _5490_ (.A1(_0778_),
    .A2(_0534_),
    .B1(_0584_),
    .B2(_0537_),
    .Y(_1894_));
 sky130_fd_sc_hd__a221oi_1 _5491_ (.A1(_0561_),
    .A2(_0527_),
    .B1(_0556_),
    .B2(_0531_),
    .C1(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__and4_1 _5492_ (.A(_1885_),
    .B(_1890_),
    .C(_1893_),
    .D(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__nand2_1 _5493_ (.A(_0554_),
    .B(_3090_),
    .Y(_1897_));
 sky130_fd_sc_hd__nand2_1 _5494_ (.A(_0559_),
    .B(_3087_),
    .Y(_1898_));
 sky130_fd_sc_hd__nand2_1 _5495_ (.A(_1897_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__a221oi_1 _5496_ (.A1(_3093_),
    .A2(_0547_),
    .B1(_3098_),
    .B2(_0551_),
    .C1(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__nand2_1 _5497_ (.A(_0573_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2_1 _5498_ (.A(_0578_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1902_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_1901_),
    .B(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__a221oi_1 _5500_ (.A1(_0542_),
    .A2(_0567_),
    .B1(_0549_),
    .B2(_0570_),
    .C1(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__nand2_1 _5501_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _5502_ (.A(_0593_),
    .B(_3072_),
    .Y(_1906_));
 sky130_fd_sc_hd__or2_1 _5503_ (.A(_0610_),
    .B(_0598_),
    .X(_1907_));
 sky130_fd_sc_hd__o2111a_1 _5504_ (.A1(_0737_),
    .A2(_0585_),
    .B1(_1905_),
    .C1(_1906_),
    .D1(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__nand2_1 _5505_ (.A(_0614_),
    .B(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1909_));
 sky130_fd_sc_hd__o21ai_1 _5506_ (.A1(_1145_),
    .A2(_0611_),
    .B1(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hd__a221oi_1 _5507_ (.A1(_3101_),
    .A2(_0604_),
    .B1(_3104_),
    .B2(_0608_),
    .C1(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__and4_1 _5508_ (.A(_1900_),
    .B(_1904_),
    .C(_1908_),
    .D(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__and4_1 _5509_ (.A(_1872_),
    .B(_1883_),
    .C(_1896_),
    .D(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__nand2_1 _5510_ (.A(_0623_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1914_));
 sky130_fd_sc_hd__nand3_1 _5511_ (.A(_1857_),
    .B(_1913_),
    .C(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__nor2_1 _5512_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__nor2_1 _5513_ (.A(_1799_),
    .B(_1916_),
    .Y(_0287_));
 sky130_fd_sc_hd__o21ai_1 _5514_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .A2(_3070_),
    .B1(_3009_),
    .Y(_1917_));
 sky130_fd_sc_hd__nand2_1 _5515_ (.A(_3153_),
    .B(_0677_),
    .Y(_1918_));
 sky130_fd_sc_hd__a22o_1 _5516_ (.A1(_3160_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .B1(_3165_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_1919_));
 sky130_fd_sc_hd__inv_2 _5517_ (.A(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__o211a_1 _5518_ (.A1(_0676_),
    .A2(_3146_),
    .B1(_1918_),
    .C1(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__nand2_1 _5519_ (.A(_3189_),
    .B(_3222_),
    .Y(_1922_));
 sky130_fd_sc_hd__o21ai_1 _5520_ (.A1(_1193_),
    .A2(_3185_),
    .B1(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__a221oi_1 _5521_ (.A1(_3167_),
    .A2(_3175_),
    .B1(_3241_),
    .B2(_3180_),
    .C1(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__nand2_1 _5522_ (.A(_3203_),
    .B(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_1925_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(_3210_),
    .B(_3227_),
    .Y(_1926_));
 sky130_fd_sc_hd__or2_1 _5524_ (.A(_1560_),
    .B(_3218_),
    .X(_1927_));
 sky130_fd_sc_hd__o2111a_1 _5525_ (.A1(_3359_),
    .A2(_3199_),
    .B1(_1925_),
    .C1(_1926_),
    .D1(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__nand2_1 _5526_ (.A(_3233_),
    .B(_3347_),
    .Y(_1929_));
 sky130_fd_sc_hd__nand2_1 _5527_ (.A(_3239_),
    .B(_3318_),
    .Y(_1930_));
 sky130_fd_sc_hd__nand2_1 _5528_ (.A(_1929_),
    .B(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__a221oi_1 _5529_ (.A1(_3342_),
    .A2(_3225_),
    .B1(_3331_),
    .B2(_3229_),
    .C1(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__and4_1 _5530_ (.A(_1921_),
    .B(_1924_),
    .C(_1928_),
    .D(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__nand2_1 _5531_ (.A(_3254_),
    .B(_3177_),
    .Y(_1934_));
 sky130_fd_sc_hd__nand2_1 _5532_ (.A(_3259_),
    .B(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_1935_));
 sky130_fd_sc_hd__or2_1 _5533_ (.A(_3183_),
    .B(_3264_),
    .X(_1936_));
 sky130_fd_sc_hd__o2111a_1 _5534_ (.A1(_0961_),
    .A2(_3251_),
    .B1(_1934_),
    .C1(_1935_),
    .D1(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__nand2_1 _5535_ (.A(_3272_),
    .B(_3214_),
    .Y(_1938_));
 sky130_fd_sc_hd__nand2_1 _5536_ (.A(_3276_),
    .B(_3191_),
    .Y(_1939_));
 sky130_fd_sc_hd__or2_1 _5537_ (.A(_0797_),
    .B(_3280_),
    .X(_1940_));
 sky130_fd_sc_hd__o2111a_1 _5538_ (.A1(_0642_),
    .A2(_3269_),
    .B1(_1938_),
    .C1(_1939_),
    .D1(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__or2_1 _5539_ (.A(_0664_),
    .B(_3293_),
    .X(_1942_));
 sky130_fd_sc_hd__o221a_1 _5540_ (.A1(_3306_),
    .A2(_3286_),
    .B1(_3303_),
    .B2(_3289_),
    .C1(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__o22ai_1 _5541_ (.A1(_3196_),
    .A2(_3304_),
    .B1(_3136_),
    .B2(_3307_),
    .Y(_1944_));
 sky130_fd_sc_hd__a221oi_1 _5542_ (.A1(_3155_),
    .A2(_3298_),
    .B1(_0631_),
    .B2(_3301_),
    .C1(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__and4_1 _5543_ (.A(_1937_),
    .B(_1941_),
    .C(_1943_),
    .D(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__o22ai_1 _5544_ (.A1(_3377_),
    .A2(_3323_),
    .B1(_3431_),
    .B2(_3327_),
    .Y(_1947_));
 sky130_fd_sc_hd__a221oi_1 _5545_ (.A1(_1107_),
    .A2(_3316_),
    .B1(_3423_),
    .B2(_3320_),
    .C1(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand2_1 _5546_ (.A(_3340_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1949_));
 sky130_fd_sc_hd__nand2_1 _5547_ (.A(_3345_),
    .B(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _5548_ (.A(_1949_),
    .B(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hd__a221oi_1 _5549_ (.A1(_0689_),
    .A2(_3333_),
    .B1(_3394_),
    .B2(_3337_),
    .C1(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__nand2_1 _5550_ (.A(_3363_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1953_));
 sky130_fd_sc_hd__o21ai_1 _5551_ (.A1(_1590_),
    .A2(_3360_),
    .B1(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__a221oi_1 _5552_ (.A1(_3335_),
    .A2(_3353_),
    .B1(_3369_),
    .B2(_3357_),
    .C1(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand2_1 _5553_ (.A(_3381_),
    .B(_0980_),
    .Y(_1956_));
 sky130_fd_sc_hd__o21ai_1 _5554_ (.A1(_0698_),
    .A2(_3378_),
    .B1(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__a221oi_1 _5555_ (.A1(_0687_),
    .A2(_3371_),
    .B1(_0839_),
    .B2(_3375_),
    .C1(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__and4_1 _5556_ (.A(_1948_),
    .B(_1952_),
    .C(_1955_),
    .D(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__nand2_1 _5557_ (.A(_3392_),
    .B(_0370_),
    .Y(_1960_));
 sky130_fd_sc_hd__nand2_1 _5558_ (.A(_3397_),
    .B(_0853_),
    .Y(_1961_));
 sky130_fd_sc_hd__or2_1 _5559_ (.A(_0863_),
    .B(_3402_),
    .X(_1962_));
 sky130_fd_sc_hd__o2111a_1 _5560_ (.A1(_0364_),
    .A2(_3389_),
    .B1(_1960_),
    .C1(_1961_),
    .D1(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__nand2_1 _5561_ (.A(_3410_),
    .B(_0360_),
    .Y(_1964_));
 sky130_fd_sc_hd__nand2_1 _5562_ (.A(_3414_),
    .B(_0718_),
    .Y(_1965_));
 sky130_fd_sc_hd__or2_1 _5563_ (.A(_1132_),
    .B(_3419_),
    .X(_1966_));
 sky130_fd_sc_hd__o2111a_1 _5564_ (.A1(_0722_),
    .A2(_3407_),
    .B1(_1964_),
    .C1(_1965_),
    .D1(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__nand2_1 _5565_ (.A(_3435_),
    .B(_3440_),
    .Y(_1968_));
 sky130_fd_sc_hd__o21ai_1 _5566_ (.A1(_3406_),
    .A2(_3432_),
    .B1(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__a221oi_1 _5567_ (.A1(_0322_),
    .A2(_3425_),
    .B1(_0705_),
    .B2(_3429_),
    .C1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _5568_ (.A(_0330_),
    .B(_0350_),
    .Y(_1971_));
 sky130_fd_sc_hd__o21ai_1 _5569_ (.A1(_0711_),
    .A2(_0327_),
    .B1(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__a221oi_1 _5570_ (.A1(_0720_),
    .A2(_3442_),
    .B1(_0868_),
    .B2(_0324_),
    .C1(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__and4_1 _5571_ (.A(_1963_),
    .B(_1967_),
    .C(_1970_),
    .D(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__and4_1 _5572_ (.A(_1933_),
    .B(_1946_),
    .C(_1959_),
    .D(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__o22ai_1 _5573_ (.A1(_1858_),
    .A2(_0348_),
    .B1(_0511_),
    .B2(_0352_),
    .Y(_1976_));
 sky130_fd_sc_hd__a221oi_1 _5574_ (.A1(_0897_),
    .A2(_0341_),
    .B1(_1032_),
    .B2(_0345_),
    .C1(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _5575_ (.A(_0368_),
    .B(_0408_),
    .Y(_1978_));
 sky130_fd_sc_hd__o21ai_1 _5576_ (.A1(_0860_),
    .A2(_0365_),
    .B1(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__a221oi_1 _5577_ (.A1(_0403_),
    .A2(_0358_),
    .B1(_0392_),
    .B2(_0362_),
    .C1(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _5578_ (.A(_0378_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1981_));
 sky130_fd_sc_hd__nand2_1 _5579_ (.A(_0383_),
    .B(_0872_),
    .Y(_1982_));
 sky130_fd_sc_hd__or2_1 _5580_ (.A(_1498_),
    .B(_0388_),
    .X(_1983_));
 sky130_fd_sc_hd__o2111a_1 _5581_ (.A1(_1740_),
    .A2(_0375_),
    .B1(_1981_),
    .C1(_1982_),
    .D1(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__nand2_1 _5582_ (.A(_0401_),
    .B(_0758_),
    .Y(_1985_));
 sky130_fd_sc_hd__nand2_1 _5583_ (.A(_0406_),
    .B(_0522_),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_1 _5584_ (.A(_1985_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__a221oi_1 _5585_ (.A1(_0904_),
    .A2(_0394_),
    .B1(_0474_),
    .B2(_0398_),
    .C1(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__and4_1 _5586_ (.A(_1977_),
    .B(_1980_),
    .C(_1984_),
    .D(_1988_),
    .X(_1989_));
 sky130_fd_sc_hd__o22ai_1 _5587_ (.A1(_0888_),
    .A2(_0422_),
    .B1(_1025_),
    .B2(_0425_),
    .Y(_1990_));
 sky130_fd_sc_hd__a221oi_1 _5588_ (.A1(_0787_),
    .A2(_0416_),
    .B1(_3284_),
    .B2(_0419_),
    .C1(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand2_1 _5589_ (.A(_0439_),
    .B(_3246_),
    .Y(_1992_));
 sky130_fd_sc_hd__o21ai_1 _5590_ (.A1(_0650_),
    .A2(_0436_),
    .B1(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__a221oi_1 _5591_ (.A1(_3291_),
    .A2(_0430_),
    .B1(_3261_),
    .B2(_0433_),
    .C1(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__nand2_1 _5592_ (.A(_0454_),
    .B(_3119_),
    .Y(_1995_));
 sky130_fd_sc_hd__o21ai_1 _5593_ (.A1(_0435_),
    .A2(_0451_),
    .B1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__a221oi_1 _5594_ (.A1(_3122_),
    .A2(_0445_),
    .B1(_3125_),
    .B2(_0448_),
    .C1(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__o22ai_1 _5595_ (.A1(_3263_),
    .A2(_0466_),
    .B1(_0653_),
    .B2(_0469_),
    .Y(_1998_));
 sky130_fd_sc_hd__a221oi_1 _5596_ (.A1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .A2(_0460_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .B2(_0463_),
    .C1(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__and4_1 _5597_ (.A(_1991_),
    .B(_1994_),
    .C(_1997_),
    .D(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__o22ai_1 _5598_ (.A1(_1412_),
    .A2(_0486_),
    .B1(_1534_),
    .B2(_0489_),
    .Y(_2001_));
 sky130_fd_sc_hd__a221oi_1 _5599_ (.A1(_0774_),
    .A2(_0479_),
    .B1(_0595_),
    .B2(_0483_),
    .C1(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__nand2_1 _5600_ (.A(_0494_),
    .B(_0745_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(_0498_),
    .B(_0525_),
    .Y(_2004_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_0503_),
    .B(_0481_),
    .Y(_2005_));
 sky130_fd_sc_hd__nand2_1 _5603_ (.A(_0507_),
    .B(_0892_),
    .Y(_2006_));
 sky130_fd_sc_hd__and4_1 _5604_ (.A(_2003_),
    .B(_2004_),
    .C(_2005_),
    .D(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__o22ai_1 _5605_ (.A1(_0907_),
    .A2(_0512_),
    .B1(_1040_),
    .B2(_0515_),
    .Y(_2008_));
 sky130_fd_sc_hd__a22o_1 _5606_ (.A1(_0518_),
    .A2(_0569_),
    .B1(_0520_),
    .B2(_0580_),
    .X(_2009_));
 sky130_fd_sc_hd__nor2_1 _5607_ (.A(_2008_),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__o22ai_1 _5608_ (.A1(_0584_),
    .A2(_0534_),
    .B1(_0773_),
    .B2(_0537_),
    .Y(_2011_));
 sky130_fd_sc_hd__a221oi_1 _5609_ (.A1(_0556_),
    .A2(_0527_),
    .B1(_0542_),
    .B2(_0531_),
    .C1(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__and4_1 _5610_ (.A(_2002_),
    .B(_2007_),
    .C(_2010_),
    .D(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__nand2_1 _5611_ (.A(_0554_),
    .B(_3093_),
    .Y(_2014_));
 sky130_fd_sc_hd__nand2_1 _5612_ (.A(_0559_),
    .B(_3090_),
    .Y(_2015_));
 sky130_fd_sc_hd__nand2_1 _5613_ (.A(_2014_),
    .B(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__a221oi_1 _5614_ (.A1(_3098_),
    .A2(_0547_),
    .B1(_3101_),
    .B2(_0551_),
    .C1(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(_0573_),
    .B(_0781_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand2_1 _5616_ (.A(_0578_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _5617_ (.A(_2018_),
    .B(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__a221oi_1 _5618_ (.A1(_0549_),
    .A2(_0567_),
    .B1(_0602_),
    .B2(_0570_),
    .C1(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_1 _5619_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_1 _5620_ (.A(_0593_),
    .B(_3084_),
    .Y(_2023_));
 sky130_fd_sc_hd__or2_1 _5621_ (.A(_0450_),
    .B(_0598_),
    .X(_2024_));
 sky130_fd_sc_hd__o2111a_1 _5622_ (.A1(_0884_),
    .A2(_0585_),
    .B1(_2022_),
    .C1(_2023_),
    .D1(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__nand2_1 _5623_ (.A(_0614_),
    .B(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_2026_));
 sky130_fd_sc_hd__o21ai_1 _5624_ (.A1(_1268_),
    .A2(_0611_),
    .B1(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__a221oi_1 _5625_ (.A1(_3104_),
    .A2(_0604_),
    .B1(_3107_),
    .B2(_0608_),
    .C1(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__and4_1 _5626_ (.A(_2017_),
    .B(_2021_),
    .C(_2025_),
    .D(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__and4_1 _5627_ (.A(_1989_),
    .B(_2000_),
    .C(_2013_),
    .D(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__nand2_1 _5628_ (.A(_0623_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_2031_));
 sky130_fd_sc_hd__nand3_1 _5629_ (.A(_1975_),
    .B(_2030_),
    .C(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__nor2_1 _5630_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(_2032_),
    .Y(_2033_));
 sky130_fd_sc_hd__nor2_1 _5631_ (.A(_1917_),
    .B(_2033_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_1 _5632_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(_3070_),
    .B1(_3009_),
    .Y(_2034_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_3153_),
    .B(_3325_),
    .Y(_2035_));
 sky130_fd_sc_hd__a22o_1 _5634_ (.A1(_3160_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .B1(_3165_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_2036_));
 sky130_fd_sc_hd__inv_2 _5635_ (.A(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__o211a_1 _5636_ (.A1(_3322_),
    .A2(_3146_),
    .B1(_2035_),
    .C1(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__nand2_1 _5637_ (.A(_3189_),
    .B(_3227_),
    .Y(_2039_));
 sky130_fd_sc_hd__o21ai_1 _5638_ (.A1(_1316_),
    .A2(_3185_),
    .B1(_2039_),
    .Y(_2040_));
 sky130_fd_sc_hd__a221oi_1 _5639_ (.A1(_3241_),
    .A2(_3175_),
    .B1(_3235_),
    .B2(_3180_),
    .C1(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__nand2_1 _5640_ (.A(_3203_),
    .B(_0675_),
    .Y(_2042_));
 sky130_fd_sc_hd__nand2_1 _5641_ (.A(_3210_),
    .B(_3351_),
    .Y(_2043_));
 sky130_fd_sc_hd__or2_1 _5642_ (.A(_1680_),
    .B(_3218_),
    .X(_2044_));
 sky130_fd_sc_hd__o2111a_1 _5643_ (.A1(_0676_),
    .A2(_3199_),
    .B1(_2042_),
    .C1(_2043_),
    .D1(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__nand2_1 _5644_ (.A(_3233_),
    .B(_3342_),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _5645_ (.A(_3239_),
    .B(_3347_),
    .Y(_2047_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_2046_),
    .B(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__a221oi_1 _5647_ (.A1(_3331_),
    .A2(_3225_),
    .B1(_3335_),
    .B2(_3229_),
    .C1(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__and4_1 _5648_ (.A(_2038_),
    .B(_2041_),
    .C(_2045_),
    .D(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__nand2_1 _5649_ (.A(_3254_),
    .B(_3182_),
    .Y(_2051_));
 sky130_fd_sc_hd__nand2_1 _5650_ (.A(_3259_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_2052_));
 sky130_fd_sc_hd__or2_1 _5651_ (.A(_0636_),
    .B(_3264_),
    .X(_2053_));
 sky130_fd_sc_hd__o2111a_1 _5652_ (.A1(_1093_),
    .A2(_3251_),
    .B1(_2051_),
    .C1(_2052_),
    .D1(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__nand2_1 _5653_ (.A(_3272_),
    .B(_3205_),
    .Y(_2055_));
 sky130_fd_sc_hd__nand2_1 _5654_ (.A(_3276_),
    .B(_3212_),
    .Y(_2056_));
 sky130_fd_sc_hd__or2_1 _5655_ (.A(_3215_),
    .B(_3280_),
    .X(_2057_));
 sky130_fd_sc_hd__o2111a_1 _5656_ (.A1(_3196_),
    .A2(_3269_),
    .B1(_2055_),
    .C1(_2056_),
    .D1(_2057_),
    .X(_2058_));
 sky130_fd_sc_hd__or2_1 _5657_ (.A(_0820_),
    .B(_3293_),
    .X(_2059_));
 sky130_fd_sc_hd__o221a_1 _5658_ (.A1(_0664_),
    .A2(_3286_),
    .B1(_3306_),
    .B2(_3289_),
    .C1(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__o22ai_1 _5659_ (.A1(_3136_),
    .A2(_3304_),
    .B1(_0630_),
    .B2(_3307_),
    .Y(_2061_));
 sky130_fd_sc_hd__a221oi_1 _5660_ (.A1(_0631_),
    .A2(_3298_),
    .B1(_3167_),
    .B2(_3301_),
    .C1(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__and4_1 _5661_ (.A(_2054_),
    .B(_2058_),
    .C(_2060_),
    .D(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__o22ai_1 _5662_ (.A1(_3431_),
    .A2(_3323_),
    .B1(_0701_),
    .B2(_3327_),
    .Y(_2064_));
 sky130_fd_sc_hd__a221oi_1 _5663_ (.A1(_3423_),
    .A2(_3316_),
    .B1(_3427_),
    .B2(_3320_),
    .C1(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__nand2_1 _5664_ (.A(_3340_),
    .B(_0689_),
    .Y(_2066_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(_3345_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_2067_));
 sky130_fd_sc_hd__nand2_1 _5666_ (.A(_2066_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__a221oi_1 _5667_ (.A1(_3394_),
    .A2(_3333_),
    .B1(_0687_),
    .B2(_3337_),
    .C1(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__nand2_1 _5668_ (.A(_3363_),
    .B(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_2070_));
 sky130_fd_sc_hd__o21ai_1 _5669_ (.A1(_1710_),
    .A2(_3360_),
    .B1(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__a221oi_1 _5670_ (.A1(_3369_),
    .A2(_3353_),
    .B1(_3373_),
    .B2(_3357_),
    .C1(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__nand2_1 _5671_ (.A(_3381_),
    .B(_3416_),
    .Y(_2073_));
 sky130_fd_sc_hd__o21ai_1 _5672_ (.A1(_3406_),
    .A2(_3378_),
    .B1(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__a221oi_1 _5673_ (.A1(_0839_),
    .A2(_3371_),
    .B1(_0980_),
    .B2(_3375_),
    .C1(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__and4_1 _5674_ (.A(_2065_),
    .B(_2069_),
    .C(_2072_),
    .D(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_3392_),
    .B(_0356_),
    .Y(_2077_));
 sky130_fd_sc_hd__nand2_1 _5676_ (.A(_3397_),
    .B(_0854_),
    .Y(_2078_));
 sky130_fd_sc_hd__or2_1 _5677_ (.A(_1002_),
    .B(_3402_),
    .X(_2079_));
 sky130_fd_sc_hd__o2111a_1 _5678_ (.A1(_0714_),
    .A2(_3389_),
    .B1(_2077_),
    .C1(_2078_),
    .D1(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__nand2_1 _5679_ (.A(_3410_),
    .B(_0380_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_1 _5680_ (.A(_3414_),
    .B(_0385_),
    .Y(_2082_));
 sky130_fd_sc_hd__or2_1 _5681_ (.A(_0387_),
    .B(_3419_),
    .X(_2083_));
 sky130_fd_sc_hd__o2111a_1 _5682_ (.A1(_0374_),
    .A2(_3407_),
    .B1(_2081_),
    .C1(_2082_),
    .D1(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__nand2_1 _5683_ (.A(_3435_),
    .B(_0322_),
    .Y(_2085_));
 sky130_fd_sc_hd__o21ai_1 _5684_ (.A1(_0694_),
    .A2(_3432_),
    .B1(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__a221oi_1 _5685_ (.A1(_0705_),
    .A2(_3425_),
    .B1(_0853_),
    .B2(_3429_),
    .C1(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__nand2_1 _5686_ (.A(_0330_),
    .B(_0337_),
    .Y(_2088_));
 sky130_fd_sc_hd__o21ai_1 _5687_ (.A1(_0860_),
    .A2(_0327_),
    .B1(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__a221oi_1 _5688_ (.A1(_0868_),
    .A2(_3442_),
    .B1(_0350_),
    .B2(_0324_),
    .C1(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__and4_1 _5689_ (.A(_2080_),
    .B(_2084_),
    .C(_2087_),
    .D(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__and4_1 _5690_ (.A(_2050_),
    .B(_2063_),
    .C(_2076_),
    .D(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__o22ai_1 _5691_ (.A1(_0511_),
    .A2(_0348_),
    .B1(_0514_),
    .B2(_0352_),
    .Y(_2093_));
 sky130_fd_sc_hd__a221oi_1 _5692_ (.A1(_1032_),
    .A2(_0341_),
    .B1(_0522_),
    .B2(_0345_),
    .C1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__nand2_1 _5693_ (.A(_0368_),
    .B(_0403_),
    .Y(_2095_));
 sky130_fd_sc_hd__o21ai_1 _5694_ (.A1(_0999_),
    .A2(_0365_),
    .B1(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__a221oi_2 _5695_ (.A1(_0392_),
    .A2(_0358_),
    .B1(_0396_),
    .B2(_0362_),
    .C1(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__nand2_1 _5696_ (.A(_0378_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_2098_));
 sky130_fd_sc_hd__nand2_1 _5697_ (.A(_0383_),
    .B(_0749_),
    .Y(_2099_));
 sky130_fd_sc_hd__or2_1 _5698_ (.A(_1620_),
    .B(_0388_),
    .X(_2100_));
 sky130_fd_sc_hd__o2111a_1 _5699_ (.A1(_1858_),
    .A2(_0375_),
    .B1(_2098_),
    .C1(_2099_),
    .D1(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__nand2_1 _5700_ (.A(_0401_),
    .B(_0904_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand2_1 _5701_ (.A(_0406_),
    .B(_0758_),
    .Y(_2103_));
 sky130_fd_sc_hd__nand2_1 _5702_ (.A(_2102_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__a221oi_1 _5703_ (.A1(_0474_),
    .A2(_0394_),
    .B1(_0481_),
    .B2(_0398_),
    .C1(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__and4_1 _5704_ (.A(_2094_),
    .B(_2097_),
    .C(_2101_),
    .D(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__o22ai_1 _5705_ (.A1(_1025_),
    .A2(_0422_),
    .B1(_3288_),
    .B2(_0425_),
    .Y(_2107_));
 sky130_fd_sc_hd__a221oi_1 _5706_ (.A1(_3284_),
    .A2(_0416_),
    .B1(_3291_),
    .B2(_0419_),
    .C1(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__nand2_1 _5707_ (.A(_0439_),
    .B(_3256_),
    .Y(_2109_));
 sky130_fd_sc_hd__o21ai_1 _5708_ (.A1(_3263_),
    .A2(_0436_),
    .B1(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__a221oi_1 _5709_ (.A1(_3261_),
    .A2(_0430_),
    .B1(_3246_),
    .B2(_0433_),
    .C1(_2110_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_1 _5710_ (.A(_0454_),
    .B(_3122_),
    .Y(_2112_));
 sky130_fd_sc_hd__o21ai_1 _5711_ (.A1(_0465_),
    .A2(_0451_),
    .B1(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__a221oi_1 _5712_ (.A1(_3125_),
    .A2(_0445_),
    .B1(_3129_),
    .B2(_0448_),
    .C1(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__o22ai_1 _5713_ (.A1(_0653_),
    .A2(_0466_),
    .B1(_3279_),
    .B2(_0469_),
    .Y(_2115_));
 sky130_fd_sc_hd__a221oi_1 _5714_ (.A1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .A2(_0460_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .B2(_0463_),
    .C1(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__and4_1 _5715_ (.A(_2108_),
    .B(_2111_),
    .C(_2114_),
    .D(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__o22ai_1 _5716_ (.A1(_1534_),
    .A2(_0486_),
    .B1(_0597_),
    .B2(_0489_),
    .Y(_2118_));
 sky130_fd_sc_hd__a221oi_1 _5717_ (.A1(_0595_),
    .A2(_0479_),
    .B1(_0776_),
    .B2(_0483_),
    .C1(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__nand2_1 _5718_ (.A(_0494_),
    .B(_0892_),
    .Y(_2120_));
 sky130_fd_sc_hd__nand2_1 _5719_ (.A(_0498_),
    .B(_0529_),
    .Y(_2121_));
 sky130_fd_sc_hd__nand2_1 _5720_ (.A(_0503_),
    .B(_0745_),
    .Y(_2122_));
 sky130_fd_sc_hd__nand2_1 _5721_ (.A(_0507_),
    .B(_0525_),
    .Y(_2123_));
 sky130_fd_sc_hd__and4_1 _5722_ (.A(_2120_),
    .B(_2121_),
    .C(_2122_),
    .D(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__o22ai_1 _5723_ (.A1(_1040_),
    .A2(_0512_),
    .B1(_1167_),
    .B2(_0515_),
    .Y(_2125_));
 sky130_fd_sc_hd__a22o_1 _5724_ (.A1(_0518_),
    .A2(_0580_),
    .B1(_0520_),
    .B2(_0575_),
    .X(_2126_));
 sky130_fd_sc_hd__nor2_1 _5725_ (.A(_2125_),
    .B(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__o22ai_1 _5726_ (.A1(_0773_),
    .A2(_0534_),
    .B1(_0919_),
    .B2(_0537_),
    .Y(_2128_));
 sky130_fd_sc_hd__a221oi_1 _5727_ (.A1(_0542_),
    .A2(_0527_),
    .B1(_0549_),
    .B2(_0531_),
    .C1(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__and4_1 _5728_ (.A(_2119_),
    .B(_2124_),
    .C(_2127_),
    .D(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_1 _5729_ (.A(_0554_),
    .B(_3098_),
    .Y(_2131_));
 sky130_fd_sc_hd__nand2_1 _5730_ (.A(_0559_),
    .B(_3093_),
    .Y(_2132_));
 sky130_fd_sc_hd__nand2_1 _5731_ (.A(_2131_),
    .B(_2132_),
    .Y(_2133_));
 sky130_fd_sc_hd__a221oi_1 _5732_ (.A1(_3101_),
    .A2(_0547_),
    .B1(_3104_),
    .B2(_0551_),
    .C1(_2133_),
    .Y(_2134_));
 sky130_fd_sc_hd__nand2_1 _5733_ (.A(_0573_),
    .B(_0924_),
    .Y(_2135_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_0578_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_2136_));
 sky130_fd_sc_hd__nand2_1 _5735_ (.A(_2135_),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__a221oi_1 _5736_ (.A1(_0602_),
    .A2(_0567_),
    .B1(_0606_),
    .B2(_0570_),
    .C1(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__nand2_1 _5737_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_2139_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_0593_),
    .B(_3087_),
    .Y(_2140_));
 sky130_fd_sc_hd__or2_1 _5739_ (.A(_0737_),
    .B(_0598_),
    .X(_2141_));
 sky130_fd_sc_hd__o2111a_1 _5740_ (.A1(_1021_),
    .A2(_0585_),
    .B1(_2139_),
    .C1(_2140_),
    .D1(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(_0614_),
    .B(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_2143_));
 sky130_fd_sc_hd__o21ai_1 _5742_ (.A1(_0435_),
    .A2(_0611_),
    .B1(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__a221oi_1 _5743_ (.A1(_3107_),
    .A2(_0604_),
    .B1(_3110_),
    .B2(_0608_),
    .C1(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__and4_1 _5744_ (.A(_2134_),
    .B(_2138_),
    .C(_2142_),
    .D(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__and4_1 _5745_ (.A(_2106_),
    .B(_2117_),
    .C(_2130_),
    .D(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__nand2_1 _5746_ (.A(_0623_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_2148_));
 sky130_fd_sc_hd__nand3_2 _5747_ (.A(_2092_),
    .B(_2147_),
    .C(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__nor2_1 _5748_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__nor2_1 _5749_ (.A(_2034_),
    .B(_2150_),
    .Y(_0285_));
 sky130_fd_sc_hd__o21ai_1 _5750_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .A2(_3070_),
    .B1(_3009_),
    .Y(_2151_));
 sky130_fd_sc_hd__nand2_1 _5751_ (.A(_3153_),
    .B(_3312_),
    .Y(_2152_));
 sky130_fd_sc_hd__a22o_1 _5752_ (.A1(_3160_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .B1(_3165_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_2153_));
 sky130_fd_sc_hd__inv_2 _5753_ (.A(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hd__o211a_1 _5754_ (.A1(_3326_),
    .A2(_3146_),
    .B1(_2152_),
    .C1(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__nand2_1 _5755_ (.A(_3189_),
    .B(_3351_),
    .Y(_2156_));
 sky130_fd_sc_hd__o21ai_1 _5756_ (.A1(_1438_),
    .A2(_3185_),
    .B1(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__a221oi_1 _5757_ (.A1(_3235_),
    .A2(_3175_),
    .B1(_3222_),
    .B2(_3180_),
    .C1(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(_3203_),
    .B(_3365_),
    .Y(_2159_));
 sky130_fd_sc_hd__nand2_1 _5759_ (.A(_3210_),
    .B(_3355_),
    .Y(_2160_));
 sky130_fd_sc_hd__or2_1 _5760_ (.A(_3359_),
    .B(_3218_),
    .X(_2161_));
 sky130_fd_sc_hd__o2111a_1 _5761_ (.A1(_3322_),
    .A2(_3199_),
    .B1(_2159_),
    .C1(_2160_),
    .D1(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__nand2_1 _5762_ (.A(_3233_),
    .B(_3331_),
    .Y(_2163_));
 sky130_fd_sc_hd__nand2_1 _5763_ (.A(_3239_),
    .B(_3342_),
    .Y(_2164_));
 sky130_fd_sc_hd__nand2_1 _5764_ (.A(_2163_),
    .B(_2164_),
    .Y(_2165_));
 sky130_fd_sc_hd__a221oi_1 _5765_ (.A1(_3335_),
    .A2(_3225_),
    .B1(_3369_),
    .B2(_3229_),
    .C1(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__and4_1 _5766_ (.A(_2155_),
    .B(_2158_),
    .C(_2162_),
    .D(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(_3254_),
    .B(_3191_),
    .Y(_2168_));
 sky130_fd_sc_hd__nand2_1 _5768_ (.A(_3259_),
    .B(_3177_),
    .Y(_2169_));
 sky130_fd_sc_hd__or2_1 _5769_ (.A(_0797_),
    .B(_3264_),
    .X(_2170_));
 sky130_fd_sc_hd__o2111a_1 _5770_ (.A1(_3183_),
    .A2(_3251_),
    .B1(_2168_),
    .C1(_2169_),
    .D1(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__nand2_1 _5771_ (.A(_3272_),
    .B(_3195_),
    .Y(_2172_));
 sky130_fd_sc_hd__nand2_1 _5772_ (.A(_3276_),
    .B(_3214_),
    .Y(_2173_));
 sky130_fd_sc_hd__or2_1 _5773_ (.A(_0642_),
    .B(_3280_),
    .X(_2174_));
 sky130_fd_sc_hd__o2111a_1 _5774_ (.A1(_3136_),
    .A2(_3269_),
    .B1(_2172_),
    .C1(_2173_),
    .D1(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__or2_1 _5775_ (.A(_0961_),
    .B(_3293_),
    .X(_2176_));
 sky130_fd_sc_hd__o221a_1 _5776_ (.A1(_0820_),
    .A2(_3286_),
    .B1(_0664_),
    .B2(_3289_),
    .C1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__o22ai_1 _5777_ (.A1(_0630_),
    .A2(_3304_),
    .B1(_0792_),
    .B2(_3307_),
    .Y(_2178_));
 sky130_fd_sc_hd__a221oi_1 _5778_ (.A1(_3167_),
    .A2(_3298_),
    .B1(_3241_),
    .B2(_3301_),
    .C1(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__and4_1 _5779_ (.A(_2171_),
    .B(_2175_),
    .C(_2177_),
    .D(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__o22ai_1 _5780_ (.A1(_0701_),
    .A2(_3323_),
    .B1(_0849_),
    .B2(_3327_),
    .Y(_2181_));
 sky130_fd_sc_hd__a221oi_1 _5781_ (.A1(_3427_),
    .A2(_3316_),
    .B1(_3399_),
    .B2(_3320_),
    .C1(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__nand2_1 _5782_ (.A(_3340_),
    .B(_3394_),
    .Y(_2183_));
 sky130_fd_sc_hd__nand2_1 _5783_ (.A(_3345_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_2184_));
 sky130_fd_sc_hd__nand2_1 _5784_ (.A(_2183_),
    .B(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__a221oi_1 _5785_ (.A1(_0687_),
    .A2(_3333_),
    .B1(_0839_),
    .B2(_3337_),
    .C1(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__nand2_1 _5786_ (.A(_3363_),
    .B(_0975_),
    .Y(_2187_));
 sky130_fd_sc_hd__o21ai_1 _5787_ (.A1(_3377_),
    .A2(_3360_),
    .B1(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hd__a221oi_1 _5788_ (.A1(_3373_),
    .A2(_3353_),
    .B1(_0681_),
    .B2(_3357_),
    .C1(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__nand2_1 _5789_ (.A(_3381_),
    .B(_0696_),
    .Y(_2190_));
 sky130_fd_sc_hd__o21ai_1 _5790_ (.A1(_0694_),
    .A2(_3378_),
    .B1(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__a221oi_1 _5791_ (.A1(_0980_),
    .A2(_3371_),
    .B1(_3416_),
    .B2(_3375_),
    .C1(_2191_),
    .Y(_2192_));
 sky130_fd_sc_hd__and4_1 _5792_ (.A(_2182_),
    .B(_2186_),
    .C(_2189_),
    .D(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__nand2_1 _5793_ (.A(_3392_),
    .B(_0360_),
    .Y(_2194_));
 sky130_fd_sc_hd__nand2_1 _5794_ (.A(_3397_),
    .B(_0370_),
    .Y(_2195_));
 sky130_fd_sc_hd__or2_1 _5795_ (.A(_1132_),
    .B(_3402_),
    .X(_2196_));
 sky130_fd_sc_hd__o2111a_1 _5796_ (.A1(_0863_),
    .A2(_3389_),
    .B1(_2194_),
    .C1(_2195_),
    .D1(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__nand2_1 _5797_ (.A(_3410_),
    .B(_0718_),
    .Y(_2198_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_3414_),
    .B(_0720_),
    .Y(_2199_));
 sky130_fd_sc_hd__or2_1 _5799_ (.A(_0722_),
    .B(_3419_),
    .X(_2200_));
 sky130_fd_sc_hd__o2111a_1 _5800_ (.A1(_0347_),
    .A2(_3407_),
    .B1(_2198_),
    .C1(_2199_),
    .D1(_2200_),
    .X(_2201_));
 sky130_fd_sc_hd__nand2_1 _5801_ (.A(_3435_),
    .B(_0705_),
    .Y(_2202_));
 sky130_fd_sc_hd__o21ai_1 _5802_ (.A1(_0844_),
    .A2(_3432_),
    .B1(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__a221oi_1 _5803_ (.A1(_0853_),
    .A2(_3425_),
    .B1(_0854_),
    .B2(_3429_),
    .C1(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__nand2_1 _5804_ (.A(_0330_),
    .B(_0343_),
    .Y(_2205_));
 sky130_fd_sc_hd__o21ai_1 _5805_ (.A1(_0999_),
    .A2(_0327_),
    .B1(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__a221oi_1 _5806_ (.A1(_0350_),
    .A2(_3442_),
    .B1(_0337_),
    .B2(_0324_),
    .C1(_2206_),
    .Y(_2207_));
 sky130_fd_sc_hd__and4_1 _5807_ (.A(_2197_),
    .B(_2201_),
    .C(_2204_),
    .D(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__and4_1 _5808_ (.A(_2167_),
    .B(_2180_),
    .C(_2193_),
    .D(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__o22ai_1 _5809_ (.A1(_0514_),
    .A2(_0348_),
    .B1(_0756_),
    .B2(_0352_),
    .Y(_2210_));
 sky130_fd_sc_hd__a221oi_1 _5810_ (.A1(_0522_),
    .A2(_0341_),
    .B1(_0758_),
    .B2(_0345_),
    .C1(_2210_),
    .Y(_2211_));
 sky130_fd_sc_hd__nand2_1 _5811_ (.A(_0368_),
    .B(_0392_),
    .Y(_2212_));
 sky130_fd_sc_hd__o21ai_1 _5812_ (.A1(_1129_),
    .A2(_0365_),
    .B1(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__a221oi_1 _5813_ (.A1(_0396_),
    .A2(_0358_),
    .B1(_0725_),
    .B2(_0362_),
    .C1(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__nand2_1 _5814_ (.A(_0378_),
    .B(_0872_),
    .Y(_2215_));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(_0383_),
    .B(_0500_),
    .Y(_2216_));
 sky130_fd_sc_hd__or2_1 _5816_ (.A(_1740_),
    .B(_0388_),
    .X(_2217_));
 sky130_fd_sc_hd__o2111a_1 _5817_ (.A1(_0511_),
    .A2(_0375_),
    .B1(_2215_),
    .C1(_2216_),
    .D1(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__nand2_1 _5818_ (.A(_0401_),
    .B(_0474_),
    .Y(_2219_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_0406_),
    .B(_0904_),
    .Y(_2220_));
 sky130_fd_sc_hd__nand2_1 _5820_ (.A(_2219_),
    .B(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hd__a221oi_1 _5821_ (.A1(_0481_),
    .A2(_0394_),
    .B1(_0745_),
    .B2(_0398_),
    .C1(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__and4_1 _5822_ (.A(_2211_),
    .B(_2214_),
    .C(_2218_),
    .D(_2222_),
    .X(_2223_));
 sky130_fd_sc_hd__o22ai_1 _5823_ (.A1(_3288_),
    .A2(_0422_),
    .B1(_3285_),
    .B2(_0425_),
    .Y(_2224_));
 sky130_fd_sc_hd__a221oi_1 _5824_ (.A1(_3291_),
    .A2(_0416_),
    .B1(_3261_),
    .B2(_0419_),
    .C1(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_0439_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_2226_));
 sky130_fd_sc_hd__o21ai_1 _5826_ (.A1(_0653_),
    .A2(_0436_),
    .B1(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a221oi_1 _5827_ (.A1(_3246_),
    .A2(_0430_),
    .B1(_3256_),
    .B2(_0433_),
    .C1(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_0454_),
    .B(_3125_),
    .Y(_2229_));
 sky130_fd_sc_hd__o21ai_1 _5829_ (.A1(_0468_),
    .A2(_0451_),
    .B1(_2229_),
    .Y(_2230_));
 sky130_fd_sc_hd__a221oi_1 _5830_ (.A1(_3129_),
    .A2(_0445_),
    .B1(_0625_),
    .B2(_0448_),
    .C1(_2230_),
    .Y(_2231_));
 sky130_fd_sc_hd__o22ai_1 _5831_ (.A1(_3279_),
    .A2(_0466_),
    .B1(_0658_),
    .B2(_0469_),
    .Y(_2232_));
 sky130_fd_sc_hd__a221oi_1 _5832_ (.A1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .A2(_0460_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .B2(_0463_),
    .C1(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__and4_1 _5833_ (.A(_2225_),
    .B(_2228_),
    .C(_2231_),
    .D(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__o22ai_1 _5834_ (.A1(_0597_),
    .A2(_0486_),
    .B1(_0778_),
    .B2(_0489_),
    .Y(_2235_));
 sky130_fd_sc_hd__a221oi_1 _5835_ (.A1(_0776_),
    .A2(_0479_),
    .B1(_0561_),
    .B2(_0483_),
    .C1(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__nand2_1 _5836_ (.A(_0494_),
    .B(_0525_),
    .Y(_2237_));
 sky130_fd_sc_hd__nand2_1 _5837_ (.A(_0498_),
    .B(_0565_),
    .Y(_2238_));
 sky130_fd_sc_hd__nand2_1 _5838_ (.A(_0503_),
    .B(_0892_),
    .Y(_2239_));
 sky130_fd_sc_hd__nand2_1 _5839_ (.A(_0507_),
    .B(_0529_),
    .Y(_2240_));
 sky130_fd_sc_hd__and4_1 _5840_ (.A(_2237_),
    .B(_2238_),
    .C(_2239_),
    .D(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__o22ai_1 _5841_ (.A1(_1167_),
    .A2(_0512_),
    .B1(_1290_),
    .B2(_0515_),
    .Y(_2242_));
 sky130_fd_sc_hd__a22o_1 _5842_ (.A1(_0518_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .B1(_0520_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_2243_));
 sky130_fd_sc_hd__nor2_1 _5843_ (.A(_2242_),
    .B(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__o22ai_1 _5844_ (.A1(_0919_),
    .A2(_0534_),
    .B1(_1052_),
    .B2(_0537_),
    .Y(_2245_));
 sky130_fd_sc_hd__a221oi_1 _5845_ (.A1(_0549_),
    .A2(_0527_),
    .B1(_0602_),
    .B2(_0531_),
    .C1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__and4_1 _5846_ (.A(_2236_),
    .B(_2241_),
    .C(_2244_),
    .D(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_0554_),
    .B(_3101_),
    .Y(_2248_));
 sky130_fd_sc_hd__nand2_1 _5848_ (.A(_0559_),
    .B(_3098_),
    .Y(_2249_));
 sky130_fd_sc_hd__nand2_1 _5849_ (.A(_2248_),
    .B(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__a221oi_1 _5850_ (.A1(_3104_),
    .A2(_0547_),
    .B1(_3107_),
    .B2(_0551_),
    .C1(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_0573_),
    .B(_3072_),
    .Y(_2252_));
 sky130_fd_sc_hd__nand2_1 _5852_ (.A(_0578_),
    .B(_0924_),
    .Y(_2253_));
 sky130_fd_sc_hd__nand2_1 _5853_ (.A(_2252_),
    .B(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__a221oi_1 _5854_ (.A1(_0606_),
    .A2(_0567_),
    .B1(_0781_),
    .B2(_0570_),
    .C1(_2254_),
    .Y(_2255_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_2256_));
 sky130_fd_sc_hd__nand2_1 _5856_ (.A(_0593_),
    .B(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_2257_));
 sky130_fd_sc_hd__or2_1 _5857_ (.A(_0884_),
    .B(_0598_),
    .X(_2258_));
 sky130_fd_sc_hd__o2111a_1 _5858_ (.A1(_0421_),
    .A2(_0585_),
    .B1(_2256_),
    .C1(_2257_),
    .D1(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__nand2_1 _5859_ (.A(_0614_),
    .B(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_2260_));
 sky130_fd_sc_hd__o21ai_1 _5860_ (.A1(_0465_),
    .A2(_0611_),
    .B1(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__a221oi_1 _5861_ (.A1(_3110_),
    .A2(_0604_),
    .B1(_3113_),
    .B2(_0608_),
    .C1(_2261_),
    .Y(_2262_));
 sky130_fd_sc_hd__and4_1 _5862_ (.A(_2251_),
    .B(_2255_),
    .C(_2259_),
    .D(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__and4_1 _5863_ (.A(_2223_),
    .B(_2234_),
    .C(_2247_),
    .D(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(_0623_),
    .B(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_2265_));
 sky130_fd_sc_hd__nand3_1 _5865_ (.A(_2209_),
    .B(_2264_),
    .C(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__nor2_1 _5866_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__nor2_1 _5867_ (.A(_2151_),
    .B(_2267_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _5868_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .A2(_3070_),
    .B1(_3009_),
    .Y(_2268_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(_3153_),
    .B(_3318_),
    .Y(_2269_));
 sky130_fd_sc_hd__a22o_1 _5870_ (.A1(_3160_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .B1(_3165_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_2270_));
 sky130_fd_sc_hd__inv_2 _5871_ (.A(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__o211a_1 _5872_ (.A1(_0668_),
    .A2(_3146_),
    .B1(_2269_),
    .C1(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(_3189_),
    .B(_3355_),
    .Y(_2273_));
 sky130_fd_sc_hd__o21ai_1 _5874_ (.A1(_1560_),
    .A2(_3185_),
    .B1(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__a221oi_1 _5875_ (.A1(_3222_),
    .A2(_3175_),
    .B1(_3227_),
    .B2(_3180_),
    .C1(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_3203_),
    .B(_0677_),
    .Y(_2276_));
 sky130_fd_sc_hd__nand2_1 _5877_ (.A(_3210_),
    .B(_0675_),
    .Y(_2277_));
 sky130_fd_sc_hd__or2_1 _5878_ (.A(_0676_),
    .B(_3218_),
    .X(_2278_));
 sky130_fd_sc_hd__o2111a_1 _5879_ (.A1(_3326_),
    .A2(_3199_),
    .B1(_2276_),
    .C1(_2277_),
    .D1(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__nand2_1 _5880_ (.A(_3233_),
    .B(_3335_),
    .Y(_2280_));
 sky130_fd_sc_hd__nand2_1 _5881_ (.A(_3239_),
    .B(_3331_),
    .Y(_2281_));
 sky130_fd_sc_hd__nand2_1 _5882_ (.A(_2280_),
    .B(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__a221oi_1 _5883_ (.A1(_3369_),
    .A2(_3225_),
    .B1(_3373_),
    .B2(_3229_),
    .C1(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__and4_1 _5884_ (.A(_2272_),
    .B(_2275_),
    .C(_2279_),
    .D(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__nand2_1 _5885_ (.A(_3254_),
    .B(_3212_),
    .Y(_2285_));
 sky130_fd_sc_hd__nand2_1 _5886_ (.A(_3259_),
    .B(_3182_),
    .Y(_2286_));
 sky130_fd_sc_hd__or2_1 _5887_ (.A(_3215_),
    .B(_3264_),
    .X(_2287_));
 sky130_fd_sc_hd__o2111a_1 _5888_ (.A1(_0636_),
    .A2(_3251_),
    .B1(_2285_),
    .C1(_2286_),
    .D1(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__nand2_1 _5889_ (.A(_3272_),
    .B(_3135_),
    .Y(_2289_));
 sky130_fd_sc_hd__nand2_1 _5890_ (.A(_3276_),
    .B(_3205_),
    .Y(_2290_));
 sky130_fd_sc_hd__or2_1 _5891_ (.A(_3196_),
    .B(_3280_),
    .X(_2291_));
 sky130_fd_sc_hd__o2111a_1 _5892_ (.A1(_0630_),
    .A2(_3269_),
    .B1(_2289_),
    .C1(_2290_),
    .D1(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__or2_1 _5893_ (.A(_1093_),
    .B(_3293_),
    .X(_2293_));
 sky130_fd_sc_hd__o221a_1 _5894_ (.A1(_0961_),
    .A2(_3286_),
    .B1(_0820_),
    .B2(_3289_),
    .C1(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__o22ai_1 _5895_ (.A1(_0792_),
    .A2(_3304_),
    .B1(_0934_),
    .B2(_3307_),
    .Y(_2295_));
 sky130_fd_sc_hd__a221oi_1 _5896_ (.A1(_3241_),
    .A2(_3298_),
    .B1(_3235_),
    .B2(_3301_),
    .C1(_2295_),
    .Y(_2296_));
 sky130_fd_sc_hd__and4_1 _5897_ (.A(_2288_),
    .B(_2292_),
    .C(_2294_),
    .D(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__o22ai_1 _5898_ (.A1(_0849_),
    .A2(_3323_),
    .B1(_0990_),
    .B2(_3327_),
    .Y(_2298_));
 sky130_fd_sc_hd__a221oi_1 _5899_ (.A1(_3399_),
    .A2(_3316_),
    .B1(_0689_),
    .B2(_3320_),
    .C1(_2298_),
    .Y(_2299_));
 sky130_fd_sc_hd__nand2_1 _5900_ (.A(_3340_),
    .B(_0687_),
    .Y(_2300_));
 sky130_fd_sc_hd__nand2_1 _5901_ (.A(_3345_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_2301_));
 sky130_fd_sc_hd__nand2_1 _5902_ (.A(_2300_),
    .B(_2301_),
    .Y(_2302_));
 sky130_fd_sc_hd__a221oi_1 _5903_ (.A1(_0839_),
    .A2(_3333_),
    .B1(_0980_),
    .B2(_3337_),
    .C1(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__nand2_1 _5904_ (.A(_3363_),
    .B(_1107_),
    .Y(_2304_));
 sky130_fd_sc_hd__o21ai_1 _5905_ (.A1(_3431_),
    .A2(_3360_),
    .B1(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__a221oi_1 _5906_ (.A1(_0681_),
    .A2(_3353_),
    .B1(_0834_),
    .B2(_3357_),
    .C1(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(_3381_),
    .B(_3440_),
    .Y(_2307_));
 sky130_fd_sc_hd__o21ai_1 _5908_ (.A1(_0844_),
    .A2(_3378_),
    .B1(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__a221oi_1 _5909_ (.A1(_3416_),
    .A2(_3371_),
    .B1(_0696_),
    .B2(_3375_),
    .C1(_2308_),
    .Y(_2309_));
 sky130_fd_sc_hd__and4_1 _5910_ (.A(_2299_),
    .B(_2303_),
    .C(_2306_),
    .D(_2309_),
    .X(_2310_));
 sky130_fd_sc_hd__nand2_1 _5911_ (.A(_3392_),
    .B(_0380_),
    .Y(_2311_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(_3397_),
    .B(_0356_),
    .Y(_2312_));
 sky130_fd_sc_hd__or2_1 _5913_ (.A(_0387_),
    .B(_3402_),
    .X(_2313_));
 sky130_fd_sc_hd__o2111a_1 _5914_ (.A1(_1002_),
    .A2(_3389_),
    .B1(_2311_),
    .C1(_2312_),
    .D1(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__nand2_1 _5915_ (.A(_3410_),
    .B(_0385_),
    .Y(_2315_));
 sky130_fd_sc_hd__nand2_1 _5916_ (.A(_3414_),
    .B(_0868_),
    .Y(_2316_));
 sky130_fd_sc_hd__or2_1 _5917_ (.A(_0374_),
    .B(_3419_),
    .X(_2317_));
 sky130_fd_sc_hd__o2111a_1 _5918_ (.A1(_0351_),
    .A2(_3407_),
    .B1(_2315_),
    .C1(_2316_),
    .D1(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_3435_),
    .B(_0853_),
    .Y(_2319_));
 sky130_fd_sc_hd__o21ai_1 _5920_ (.A1(_0985_),
    .A2(_3432_),
    .B1(_2319_),
    .Y(_2320_));
 sky130_fd_sc_hd__a221oi_1 _5921_ (.A1(_0854_),
    .A2(_3425_),
    .B1(_0370_),
    .B2(_3429_),
    .C1(_2320_),
    .Y(_2321_));
 sky130_fd_sc_hd__nand2_1 _5922_ (.A(_0330_),
    .B(_0408_),
    .Y(_2322_));
 sky130_fd_sc_hd__o21ai_1 _5923_ (.A1(_1129_),
    .A2(_0327_),
    .B1(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__a221oi_1 _5924_ (.A1(_0337_),
    .A2(_3442_),
    .B1(_0343_),
    .B2(_0324_),
    .C1(_2323_),
    .Y(_2324_));
 sky130_fd_sc_hd__and4_1 _5925_ (.A(_2314_),
    .B(_2318_),
    .C(_2321_),
    .D(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__and4_1 _5926_ (.A(_2284_),
    .B(_2297_),
    .C(_2310_),
    .D(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__o22ai_1 _5927_ (.A1(_0756_),
    .A2(_0348_),
    .B1(_0902_),
    .B2(_0352_),
    .Y(_2327_));
 sky130_fd_sc_hd__a221oi_1 _5928_ (.A1(_0758_),
    .A2(_0341_),
    .B1(_0904_),
    .B2(_0345_),
    .C1(_2327_),
    .Y(_2328_));
 sky130_fd_sc_hd__nand2_1 _5929_ (.A(_0368_),
    .B(_0396_),
    .Y(_2329_));
 sky130_fd_sc_hd__o21ai_1 _5930_ (.A1(_1253_),
    .A2(_0365_),
    .B1(_2329_),
    .Y(_2330_));
 sky130_fd_sc_hd__a221oi_1 _5931_ (.A1(_0725_),
    .A2(_0358_),
    .B1(_0872_),
    .B2(_0362_),
    .C1(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__nand2_1 _5932_ (.A(_0378_),
    .B(_0749_),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _5933_ (.A(_0383_),
    .B(_0751_),
    .Y(_2333_));
 sky130_fd_sc_hd__or2_1 _5934_ (.A(_1858_),
    .B(_0388_),
    .X(_2334_));
 sky130_fd_sc_hd__o2111a_1 _5935_ (.A1(_0514_),
    .A2(_0375_),
    .B1(_2332_),
    .C1(_2333_),
    .D1(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__nand2_1 _5936_ (.A(_0401_),
    .B(_0481_),
    .Y(_2336_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(_0406_),
    .B(_0474_),
    .Y(_2337_));
 sky130_fd_sc_hd__nand2_1 _5938_ (.A(_2336_),
    .B(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__a221oi_1 _5939_ (.A1(_0745_),
    .A2(_0394_),
    .B1(_0892_),
    .B2(_0398_),
    .C1(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__and4_1 _5940_ (.A(_2328_),
    .B(_2331_),
    .C(_2335_),
    .D(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__o22ai_1 _5941_ (.A1(_3285_),
    .A2(_0422_),
    .B1(_3292_),
    .B2(_0425_),
    .Y(_2341_));
 sky130_fd_sc_hd__a221oi_1 _5942_ (.A1(_3261_),
    .A2(_0416_),
    .B1(_3246_),
    .B2(_0419_),
    .C1(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__nand2_1 _5943_ (.A(_0439_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_2343_));
 sky130_fd_sc_hd__o21ai_1 _5944_ (.A1(_3279_),
    .A2(_0436_),
    .B1(_2343_),
    .Y(_2344_));
 sky130_fd_sc_hd__a221oi_1 _5945_ (.A1(_3256_),
    .A2(_0430_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .B2(_0433_),
    .C1(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(_0454_),
    .B(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_2346_));
 sky130_fd_sc_hd__o21ai_1 _5947_ (.A1(_0741_),
    .A2(_0451_),
    .B1(_2346_),
    .Y(_2347_));
 sky130_fd_sc_hd__a221oi_1 _5948_ (.A1(_0625_),
    .A2(_0445_),
    .B1(_0787_),
    .B2(_0448_),
    .C1(_2347_),
    .Y(_2348_));
 sky130_fd_sc_hd__o22ai_1 _5949_ (.A1(_0658_),
    .A2(_0466_),
    .B1(_3268_),
    .B2(_0469_),
    .Y(_2349_));
 sky130_fd_sc_hd__a221oi_1 _5950_ (.A1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .A2(_0460_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .B2(_0463_),
    .C1(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__and4_1 _5951_ (.A(_2342_),
    .B(_2345_),
    .C(_2348_),
    .D(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__o22ai_1 _5952_ (.A1(_0778_),
    .A2(_0486_),
    .B1(_0584_),
    .B2(_0489_),
    .Y(_2352_));
 sky130_fd_sc_hd__a221oi_1 _5953_ (.A1(_0561_),
    .A2(_0479_),
    .B1(_0556_),
    .B2(_0483_),
    .C1(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__nand2_1 _5954_ (.A(_0494_),
    .B(_0529_),
    .Y(_2354_));
 sky130_fd_sc_hd__nand2_1 _5955_ (.A(_0498_),
    .B(_0569_),
    .Y(_2355_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_0503_),
    .B(_0525_),
    .Y(_2356_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(_0507_),
    .B(_0565_),
    .Y(_2357_));
 sky130_fd_sc_hd__and4_1 _5958_ (.A(_2354_),
    .B(_2355_),
    .C(_2356_),
    .D(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__o22ai_1 _5959_ (.A1(_1290_),
    .A2(_0512_),
    .B1(_1412_),
    .B2(_0515_),
    .Y(_2359_));
 sky130_fd_sc_hd__a22o_1 _5960_ (.A1(_0518_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .B1(_0520_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_2360_));
 sky130_fd_sc_hd__nor2_1 _5961_ (.A(_2359_),
    .B(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__o22ai_1 _5962_ (.A1(_1052_),
    .A2(_0534_),
    .B1(_1179_),
    .B2(_0537_),
    .Y(_2362_));
 sky130_fd_sc_hd__a221oi_1 _5963_ (.A1(_0602_),
    .A2(_0527_),
    .B1(_0606_),
    .B2(_0531_),
    .C1(_2362_),
    .Y(_2363_));
 sky130_fd_sc_hd__and4_1 _5964_ (.A(_2353_),
    .B(_2358_),
    .C(_2361_),
    .D(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_0554_),
    .B(_3104_),
    .Y(_2365_));
 sky130_fd_sc_hd__nand2_1 _5966_ (.A(_0559_),
    .B(_3101_),
    .Y(_2366_));
 sky130_fd_sc_hd__nand2_1 _5967_ (.A(_2365_),
    .B(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__a221oi_1 _5968_ (.A1(_3107_),
    .A2(_0547_),
    .B1(_3110_),
    .B2(_0551_),
    .C1(_2367_),
    .Y(_2368_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(_0573_),
    .B(_3084_),
    .Y(_2369_));
 sky130_fd_sc_hd__nand2_1 _5970_ (.A(_0578_),
    .B(_3072_),
    .Y(_2370_));
 sky130_fd_sc_hd__nand2_1 _5971_ (.A(_2369_),
    .B(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__a221oi_1 _5972_ (.A1(_0781_),
    .A2(_0567_),
    .B1(_0924_),
    .B2(_0570_),
    .C1(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__nand2_1 _5973_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_2373_));
 sky130_fd_sc_hd__nand2_1 _5974_ (.A(_0593_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_2374_));
 sky130_fd_sc_hd__or2_1 _5975_ (.A(_1021_),
    .B(_0598_),
    .X(_2375_));
 sky130_fd_sc_hd__o2111a_1 _5976_ (.A1(_0424_),
    .A2(_0585_),
    .B1(_2373_),
    .C1(_2374_),
    .D1(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__nand2_1 _5977_ (.A(_0614_),
    .B(_3119_),
    .Y(_2377_));
 sky130_fd_sc_hd__o21ai_1 _5978_ (.A1(_0468_),
    .A2(_0611_),
    .B1(_2377_),
    .Y(_2378_));
 sky130_fd_sc_hd__a221oi_1 _5979_ (.A1(_3113_),
    .A2(_0604_),
    .B1(_3116_),
    .B2(_0608_),
    .C1(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__and4_1 _5980_ (.A(_2368_),
    .B(_2372_),
    .C(_2376_),
    .D(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__and4_1 _5981_ (.A(_2340_),
    .B(_2351_),
    .C(_2364_),
    .D(_2380_),
    .X(_2381_));
 sky130_fd_sc_hd__nand2_1 _5982_ (.A(_0623_),
    .B(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_2382_));
 sky130_fd_sc_hd__nand3_2 _5983_ (.A(_2326_),
    .B(_2381_),
    .C(_2382_),
    .Y(_2383_));
 sky130_fd_sc_hd__nor2_1 _5984_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(_2383_),
    .Y(_2384_));
 sky130_fd_sc_hd__nor2_1 _5985_ (.A(_2268_),
    .B(_2384_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _5986_ (.A(_3078_),
    .B(_3052_),
    .Y(_2385_));
 sky130_fd_sc_hd__and3_1 _5987_ (.A(_3081_),
    .B(_3008_),
    .C(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__clkbuf_1 _5988_ (.A(_2386_),
    .X(_0282_));
 sky130_fd_sc_hd__nand2_1 _5989_ (.A(_3077_),
    .B(_3045_),
    .Y(_2387_));
 sky130_fd_sc_hd__and3_1 _5990_ (.A(_3078_),
    .B(_3008_),
    .C(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__clkbuf_1 _5991_ (.A(_2388_),
    .X(_0281_));
 sky130_fd_sc_hd__or2_1 _5992_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .B(_3076_),
    .X(_2389_));
 sky130_fd_sc_hd__and3_1 _5993_ (.A(_2389_),
    .B(_3008_),
    .C(_3077_),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_1 _5994_ (.A(_2390_),
    .X(_0280_));
 sky130_fd_sc_hd__nand2_4 _5995_ (.A(_3076_),
    .B(_3053_),
    .Y(_2391_));
 sky130_fd_sc_hd__clkbuf_4 _5996_ (.A(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _5997_ (.A0(net7),
    .A1(_0625_),
    .S(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__and2_1 _5998_ (.A(_2393_),
    .B(_3127_),
    .X(_2394_));
 sky130_fd_sc_hd__clkbuf_1 _5999_ (.A(_2394_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _6000_ (.A0(net6),
    .A1(_0787_),
    .S(_2392_),
    .X(_2395_));
 sky130_fd_sc_hd__and2_1 _6001_ (.A(_2395_),
    .B(_3127_),
    .X(_2396_));
 sky130_fd_sc_hd__clkbuf_1 _6002_ (.A(_2396_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _6003_ (.A0(net5),
    .A1(_3284_),
    .S(_2392_),
    .X(_2397_));
 sky130_fd_sc_hd__and2_1 _6004_ (.A(_2397_),
    .B(_3127_),
    .X(_2398_));
 sky130_fd_sc_hd__clkbuf_1 _6005_ (.A(_2398_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _6006_ (.A0(net4),
    .A1(_3291_),
    .S(_2392_),
    .X(_2399_));
 sky130_fd_sc_hd__and2_1 _6007_ (.A(_2399_),
    .B(_3127_),
    .X(_2400_));
 sky130_fd_sc_hd__clkbuf_1 _6008_ (.A(_2400_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _6009_ (.A0(net3),
    .A1(_3261_),
    .S(_2392_),
    .X(_2401_));
 sky130_fd_sc_hd__and2_1 _6010_ (.A(_2401_),
    .B(_3127_),
    .X(_2402_));
 sky130_fd_sc_hd__clkbuf_1 _6011_ (.A(_2402_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _6012_ (.A0(net2),
    .A1(_3246_),
    .S(_2392_),
    .X(_2403_));
 sky130_fd_sc_hd__and2_1 _6013_ (.A(_2403_),
    .B(_3127_),
    .X(_2404_));
 sky130_fd_sc_hd__clkbuf_1 _6014_ (.A(_2404_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _6015_ (.A0(net16),
    .A1(_3256_),
    .S(_2392_),
    .X(_2405_));
 sky130_fd_sc_hd__and2_1 _6016_ (.A(_2405_),
    .B(_3127_),
    .X(_2406_));
 sky130_fd_sc_hd__clkbuf_1 _6017_ (.A(_2406_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _6018_ (.A0(net15),
    .A1(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .S(_2392_),
    .X(_2407_));
 sky130_fd_sc_hd__and2_1 _6019_ (.A(_2407_),
    .B(_3127_),
    .X(_2408_));
 sky130_fd_sc_hd__clkbuf_1 _6020_ (.A(_2408_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _6021_ (.A0(net14),
    .A1(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .S(_2392_),
    .X(_2409_));
 sky130_fd_sc_hd__clkbuf_2 _6022_ (.A(_3095_),
    .X(_2410_));
 sky130_fd_sc_hd__and2_1 _6023_ (.A(_2409_),
    .B(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__clkbuf_1 _6024_ (.A(_2411_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _6025_ (.A0(net13),
    .A1(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .S(_2392_),
    .X(_2412_));
 sky130_fd_sc_hd__and2_1 _6026_ (.A(_2412_),
    .B(_2410_),
    .X(_2413_));
 sky130_fd_sc_hd__clkbuf_1 _6027_ (.A(_2413_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _6028_ (.A0(net12),
    .A1(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .S(_2391_),
    .X(_2414_));
 sky130_fd_sc_hd__and2_1 _6029_ (.A(_2414_),
    .B(_2410_),
    .X(_2415_));
 sky130_fd_sc_hd__clkbuf_1 _6030_ (.A(_2415_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _6031_ (.A0(net11),
    .A1(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .S(_2391_),
    .X(_2416_));
 sky130_fd_sc_hd__and2_1 _6032_ (.A(_2416_),
    .B(_2410_),
    .X(_2417_));
 sky130_fd_sc_hd__clkbuf_1 _6033_ (.A(_2417_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(net10),
    .A1(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .S(_2391_),
    .X(_2418_));
 sky130_fd_sc_hd__and2_1 _6035_ (.A(_2418_),
    .B(_2410_),
    .X(_2419_));
 sky130_fd_sc_hd__clkbuf_1 _6036_ (.A(_2419_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _6037_ (.A0(net9),
    .A1(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .S(_2391_),
    .X(_2420_));
 sky130_fd_sc_hd__and2_1 _6038_ (.A(_2420_),
    .B(_2410_),
    .X(_2421_));
 sky130_fd_sc_hd__clkbuf_1 _6039_ (.A(_2421_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _6040_ (.A0(net8),
    .A1(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .S(_2391_),
    .X(_2422_));
 sky130_fd_sc_hd__and2_1 _6041_ (.A(_2422_),
    .B(_2410_),
    .X(_2423_));
 sky130_fd_sc_hd__clkbuf_1 _6042_ (.A(_2423_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _6043_ (.A0(net1),
    .A1(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .S(_2391_),
    .X(_2424_));
 sky130_fd_sc_hd__and2_1 _6044_ (.A(_2424_),
    .B(_2410_),
    .X(_2425_));
 sky130_fd_sc_hd__clkbuf_1 _6045_ (.A(_2425_),
    .X(_0264_));
 sky130_fd_sc_hd__or4b_2 _6046_ (.A(net37),
    .B(net39),
    .C(_3046_),
    .D_N(_3076_),
    .X(_2426_));
 sky130_fd_sc_hd__buf_2 _6047_ (.A(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__clkbuf_4 _6048_ (.A(_2427_),
    .X(_2428_));
 sky130_fd_sc_hd__mux2_1 _6049_ (.A0(net7),
    .A1(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .S(_2428_),
    .X(_2429_));
 sky130_fd_sc_hd__and2_1 _6050_ (.A(_2429_),
    .B(_2410_),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_1 _6051_ (.A(_2430_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _6052_ (.A0(net6),
    .A1(_3177_),
    .S(_2428_),
    .X(_2431_));
 sky130_fd_sc_hd__and2_1 _6053_ (.A(_2431_),
    .B(_2410_),
    .X(_2432_));
 sky130_fd_sc_hd__clkbuf_1 _6054_ (.A(_2432_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _6055_ (.A0(net5),
    .A1(_3182_),
    .S(_2428_),
    .X(_2433_));
 sky130_fd_sc_hd__clkbuf_2 _6056_ (.A(_3095_),
    .X(_2434_));
 sky130_fd_sc_hd__and2_1 _6057_ (.A(_2433_),
    .B(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__clkbuf_1 _6058_ (.A(_2435_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _6059_ (.A0(net4),
    .A1(_3191_),
    .S(_2428_),
    .X(_2436_));
 sky130_fd_sc_hd__and2_1 _6060_ (.A(_2436_),
    .B(_2434_),
    .X(_2437_));
 sky130_fd_sc_hd__clkbuf_1 _6061_ (.A(_2437_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _6062_ (.A0(net3),
    .A1(_3212_),
    .S(_2428_),
    .X(_2438_));
 sky130_fd_sc_hd__and2_1 _6063_ (.A(_2438_),
    .B(_2434_),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_1 _6064_ (.A(_2439_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _6065_ (.A0(net2),
    .A1(_3214_),
    .S(_2428_),
    .X(_2440_));
 sky130_fd_sc_hd__and2_1 _6066_ (.A(_2440_),
    .B(_2434_),
    .X(_2441_));
 sky130_fd_sc_hd__clkbuf_1 _6067_ (.A(_2441_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _6068_ (.A0(net16),
    .A1(_3205_),
    .S(_2428_),
    .X(_2442_));
 sky130_fd_sc_hd__and2_1 _6069_ (.A(_2442_),
    .B(_2434_),
    .X(_2443_));
 sky130_fd_sc_hd__clkbuf_1 _6070_ (.A(_2443_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _6071_ (.A0(net15),
    .A1(_3195_),
    .S(_2428_),
    .X(_2444_));
 sky130_fd_sc_hd__and2_1 _6072_ (.A(_2444_),
    .B(_2434_),
    .X(_2445_));
 sky130_fd_sc_hd__clkbuf_1 _6073_ (.A(_2445_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _6074_ (.A0(net14),
    .A1(_3135_),
    .S(_2428_),
    .X(_2446_));
 sky130_fd_sc_hd__and2_1 _6075_ (.A(_2446_),
    .B(_2434_),
    .X(_2447_));
 sky130_fd_sc_hd__clkbuf_1 _6076_ (.A(_2447_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _6077_ (.A0(net13),
    .A1(_3155_),
    .S(_2428_),
    .X(_2448_));
 sky130_fd_sc_hd__and2_1 _6078_ (.A(_2448_),
    .B(_2434_),
    .X(_2449_));
 sky130_fd_sc_hd__clkbuf_1 _6079_ (.A(_2449_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _6080_ (.A0(net12),
    .A1(_0631_),
    .S(_2427_),
    .X(_2450_));
 sky130_fd_sc_hd__and2_1 _6081_ (.A(_2450_),
    .B(_2434_),
    .X(_2451_));
 sky130_fd_sc_hd__clkbuf_1 _6082_ (.A(_2451_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _6083_ (.A0(net11),
    .A1(_3167_),
    .S(_2427_),
    .X(_2452_));
 sky130_fd_sc_hd__and2_1 _6084_ (.A(_2452_),
    .B(_2434_),
    .X(_2453_));
 sky130_fd_sc_hd__clkbuf_1 _6085_ (.A(_2453_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _6086_ (.A0(net10),
    .A1(_3241_),
    .S(_2427_),
    .X(_2454_));
 sky130_fd_sc_hd__clkbuf_2 _6087_ (.A(_3095_),
    .X(_2455_));
 sky130_fd_sc_hd__and2_1 _6088_ (.A(_2454_),
    .B(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__clkbuf_1 _6089_ (.A(_2456_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _6090_ (.A0(net9),
    .A1(_3235_),
    .S(_2427_),
    .X(_2457_));
 sky130_fd_sc_hd__and2_1 _6091_ (.A(_2457_),
    .B(_2455_),
    .X(_2458_));
 sky130_fd_sc_hd__clkbuf_1 _6092_ (.A(_2458_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _6093_ (.A0(net8),
    .A1(_3222_),
    .S(_2427_),
    .X(_2459_));
 sky130_fd_sc_hd__and2_1 _6094_ (.A(_2459_),
    .B(_2455_),
    .X(_2460_));
 sky130_fd_sc_hd__clkbuf_1 _6095_ (.A(_2460_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _6096_ (.A0(net1),
    .A1(_3227_),
    .S(_2427_),
    .X(_2461_));
 sky130_fd_sc_hd__and2_1 _6097_ (.A(_2461_),
    .B(_2455_),
    .X(_2462_));
 sky130_fd_sc_hd__clkbuf_1 _6098_ (.A(_2462_),
    .X(_0248_));
 sky130_fd_sc_hd__or4b_2 _6099_ (.A(net37),
    .B(_3045_),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .D_N(_3076_),
    .X(_2463_));
 sky130_fd_sc_hd__buf_2 _6100_ (.A(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__clkbuf_4 _6101_ (.A(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(net7),
    .A1(_3351_),
    .S(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__and2_1 _6103_ (.A(_2466_),
    .B(_2455_),
    .X(_2467_));
 sky130_fd_sc_hd__clkbuf_1 _6104_ (.A(_2467_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _6105_ (.A0(net6),
    .A1(_3355_),
    .S(_2465_),
    .X(_2468_));
 sky130_fd_sc_hd__and2_1 _6106_ (.A(_2468_),
    .B(_2455_),
    .X(_2469_));
 sky130_fd_sc_hd__clkbuf_1 _6107_ (.A(_2469_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _6108_ (.A0(net5),
    .A1(_0675_),
    .S(_2465_),
    .X(_2470_));
 sky130_fd_sc_hd__and2_1 _6109_ (.A(_2470_),
    .B(_2455_),
    .X(_2471_));
 sky130_fd_sc_hd__clkbuf_1 _6110_ (.A(_2471_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _6111_ (.A0(net4),
    .A1(_3365_),
    .S(_2465_),
    .X(_2472_));
 sky130_fd_sc_hd__and2_1 _6112_ (.A(_2472_),
    .B(_2455_),
    .X(_2473_));
 sky130_fd_sc_hd__clkbuf_1 _6113_ (.A(_2473_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _6114_ (.A0(net3),
    .A1(_0677_),
    .S(_2465_),
    .X(_2474_));
 sky130_fd_sc_hd__and2_1 _6115_ (.A(_2474_),
    .B(_2455_),
    .X(_2475_));
 sky130_fd_sc_hd__clkbuf_1 _6116_ (.A(_2475_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _6117_ (.A0(net2),
    .A1(_3325_),
    .S(_2465_),
    .X(_2476_));
 sky130_fd_sc_hd__and2_1 _6118_ (.A(_2476_),
    .B(_2455_),
    .X(_2477_));
 sky130_fd_sc_hd__clkbuf_1 _6119_ (.A(_2477_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _6120_ (.A0(net16),
    .A1(_3312_),
    .S(_2465_),
    .X(_2478_));
 sky130_fd_sc_hd__clkbuf_2 _6121_ (.A(_3095_),
    .X(_2479_));
 sky130_fd_sc_hd__and2_1 _6122_ (.A(_2478_),
    .B(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__clkbuf_1 _6123_ (.A(_2480_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(net15),
    .A1(_3318_),
    .S(_2465_),
    .X(_2481_));
 sky130_fd_sc_hd__and2_1 _6125_ (.A(_2481_),
    .B(_2479_),
    .X(_2482_));
 sky130_fd_sc_hd__clkbuf_1 _6126_ (.A(_2482_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _6127_ (.A0(net14),
    .A1(_3347_),
    .S(_2465_),
    .X(_2483_));
 sky130_fd_sc_hd__and2_1 _6128_ (.A(_2483_),
    .B(_2479_),
    .X(_2484_));
 sky130_fd_sc_hd__clkbuf_1 _6129_ (.A(_2484_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _6130_ (.A0(net13),
    .A1(_3342_),
    .S(_2465_),
    .X(_2485_));
 sky130_fd_sc_hd__and2_1 _6131_ (.A(_2485_),
    .B(_2479_),
    .X(_2486_));
 sky130_fd_sc_hd__clkbuf_1 _6132_ (.A(_2486_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _6133_ (.A0(net12),
    .A1(_3331_),
    .S(_2464_),
    .X(_2487_));
 sky130_fd_sc_hd__and2_1 _6134_ (.A(_2487_),
    .B(_2479_),
    .X(_2488_));
 sky130_fd_sc_hd__clkbuf_1 _6135_ (.A(_2488_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _6136_ (.A0(net11),
    .A1(_3335_),
    .S(_2464_),
    .X(_2489_));
 sky130_fd_sc_hd__and2_1 _6137_ (.A(_2489_),
    .B(_2479_),
    .X(_2490_));
 sky130_fd_sc_hd__clkbuf_1 _6138_ (.A(_2490_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _6139_ (.A0(net10),
    .A1(_3369_),
    .S(_2464_),
    .X(_2491_));
 sky130_fd_sc_hd__and2_1 _6140_ (.A(_2491_),
    .B(_2479_),
    .X(_2492_));
 sky130_fd_sc_hd__clkbuf_1 _6141_ (.A(_2492_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _6142_ (.A0(net9),
    .A1(_3373_),
    .S(_2464_),
    .X(_2493_));
 sky130_fd_sc_hd__and2_1 _6143_ (.A(_2493_),
    .B(_2479_),
    .X(_2494_));
 sky130_fd_sc_hd__clkbuf_1 _6144_ (.A(_2494_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _6145_ (.A0(net8),
    .A1(_0681_),
    .S(_2464_),
    .X(_2495_));
 sky130_fd_sc_hd__and2_1 _6146_ (.A(_2495_),
    .B(_2479_),
    .X(_2496_));
 sky130_fd_sc_hd__clkbuf_1 _6147_ (.A(_2496_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _6148_ (.A0(net1),
    .A1(_0834_),
    .S(_2464_),
    .X(_2497_));
 sky130_fd_sc_hd__and2_1 _6149_ (.A(_2497_),
    .B(_2479_),
    .X(_2498_));
 sky130_fd_sc_hd__clkbuf_1 _6150_ (.A(_2498_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_2 _6151_ (.A(net37),
    .B(_3078_),
    .X(_2499_));
 sky130_fd_sc_hd__buf_2 _6152_ (.A(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__clkbuf_4 _6153_ (.A(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__mux2_1 _6154_ (.A0(net7),
    .A1(_0975_),
    .S(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__clkbuf_2 _6155_ (.A(_3095_),
    .X(_2503_));
 sky130_fd_sc_hd__and2_1 _6156_ (.A(_2502_),
    .B(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__clkbuf_1 _6157_ (.A(_2504_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _6158_ (.A0(net6),
    .A1(_1107_),
    .S(_2501_),
    .X(_2505_));
 sky130_fd_sc_hd__and2_1 _6159_ (.A(_2505_),
    .B(_2503_),
    .X(_2506_));
 sky130_fd_sc_hd__clkbuf_1 _6160_ (.A(_2506_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _6161_ (.A0(net5),
    .A1(_3423_),
    .S(_2501_),
    .X(_2507_));
 sky130_fd_sc_hd__and2_1 _6162_ (.A(_2507_),
    .B(_2503_),
    .X(_2508_));
 sky130_fd_sc_hd__clkbuf_1 _6163_ (.A(_2508_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _6164_ (.A0(net4),
    .A1(_3427_),
    .S(_2501_),
    .X(_2509_));
 sky130_fd_sc_hd__and2_1 _6165_ (.A(_2509_),
    .B(_2503_),
    .X(_2510_));
 sky130_fd_sc_hd__clkbuf_1 _6166_ (.A(_2510_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _6167_ (.A0(net3),
    .A1(_3399_),
    .S(_2501_),
    .X(_2511_));
 sky130_fd_sc_hd__and2_1 _6168_ (.A(_2511_),
    .B(_2503_),
    .X(_2512_));
 sky130_fd_sc_hd__clkbuf_1 _6169_ (.A(_2512_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _6170_ (.A0(net2),
    .A1(_0689_),
    .S(_2501_),
    .X(_2513_));
 sky130_fd_sc_hd__and2_1 _6171_ (.A(_2513_),
    .B(_2503_),
    .X(_2514_));
 sky130_fd_sc_hd__clkbuf_1 _6172_ (.A(_2514_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _6173_ (.A0(net16),
    .A1(_3394_),
    .S(_2501_),
    .X(_2515_));
 sky130_fd_sc_hd__and2_1 _6174_ (.A(_2515_),
    .B(_2503_),
    .X(_2516_));
 sky130_fd_sc_hd__clkbuf_1 _6175_ (.A(_2516_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _6176_ (.A0(net15),
    .A1(_0687_),
    .S(_2501_),
    .X(_2517_));
 sky130_fd_sc_hd__and2_1 _6177_ (.A(_2517_),
    .B(_2503_),
    .X(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _6178_ (.A(_2518_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _6179_ (.A0(net14),
    .A1(_0839_),
    .S(_2501_),
    .X(_2519_));
 sky130_fd_sc_hd__and2_1 _6180_ (.A(_2519_),
    .B(_2503_),
    .X(_2520_));
 sky130_fd_sc_hd__clkbuf_1 _6181_ (.A(_2520_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _6182_ (.A0(net13),
    .A1(_0980_),
    .S(_2501_),
    .X(_2521_));
 sky130_fd_sc_hd__and2_1 _6183_ (.A(_2521_),
    .B(_2503_),
    .X(_2522_));
 sky130_fd_sc_hd__clkbuf_1 _6184_ (.A(_2522_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _6185_ (.A0(net12),
    .A1(_3416_),
    .S(_2500_),
    .X(_2523_));
 sky130_fd_sc_hd__clkbuf_2 _6186_ (.A(_3095_),
    .X(_2524_));
 sky130_fd_sc_hd__and2_1 _6187_ (.A(_2523_),
    .B(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__clkbuf_1 _6188_ (.A(_2525_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _6189_ (.A0(net11),
    .A1(_0696_),
    .S(_2500_),
    .X(_2526_));
 sky130_fd_sc_hd__and2_1 _6190_ (.A(_2526_),
    .B(_2524_),
    .X(_2527_));
 sky130_fd_sc_hd__clkbuf_1 _6191_ (.A(_2527_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _6192_ (.A0(net10),
    .A1(_3440_),
    .S(_2500_),
    .X(_2528_));
 sky130_fd_sc_hd__and2_1 _6193_ (.A(_2528_),
    .B(_2524_),
    .X(_2529_));
 sky130_fd_sc_hd__clkbuf_1 _6194_ (.A(_2529_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _6195_ (.A0(net9),
    .A1(_0322_),
    .S(_2500_),
    .X(_2530_));
 sky130_fd_sc_hd__and2_1 _6196_ (.A(_2530_),
    .B(_2524_),
    .X(_2531_));
 sky130_fd_sc_hd__clkbuf_1 _6197_ (.A(_2531_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _6198_ (.A0(net8),
    .A1(_0705_),
    .S(_2500_),
    .X(_2532_));
 sky130_fd_sc_hd__and2_1 _6199_ (.A(_2532_),
    .B(_2524_),
    .X(_2533_));
 sky130_fd_sc_hd__clkbuf_1 _6200_ (.A(_2533_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _6201_ (.A0(net1),
    .A1(_0853_),
    .S(_2500_),
    .X(_2534_));
 sky130_fd_sc_hd__and2_1 _6202_ (.A(_2534_),
    .B(_2524_),
    .X(_2535_));
 sky130_fd_sc_hd__clkbuf_1 _6203_ (.A(_2535_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_4 _6204_ (.A(_3076_),
    .B(net38),
    .Y(_2536_));
 sky130_fd_sc_hd__clkbuf_4 _6205_ (.A(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__mux2_1 _6206_ (.A0(net7),
    .A1(_0854_),
    .S(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__and2_1 _6207_ (.A(_2538_),
    .B(_2524_),
    .X(_2539_));
 sky130_fd_sc_hd__clkbuf_1 _6208_ (.A(_2539_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _6209_ (.A0(net6),
    .A1(_0370_),
    .S(_2537_),
    .X(_2540_));
 sky130_fd_sc_hd__and2_1 _6210_ (.A(_2540_),
    .B(_2524_),
    .X(_2541_));
 sky130_fd_sc_hd__clkbuf_1 _6211_ (.A(_2541_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _6212_ (.A0(net5),
    .A1(_0356_),
    .S(_2537_),
    .X(_2542_));
 sky130_fd_sc_hd__and2_1 _6213_ (.A(_2542_),
    .B(_2524_),
    .X(_2543_));
 sky130_fd_sc_hd__clkbuf_1 _6214_ (.A(_2543_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _6215_ (.A0(net4),
    .A1(_0360_),
    .S(_2537_),
    .X(_2544_));
 sky130_fd_sc_hd__and2_1 _6216_ (.A(_2544_),
    .B(_2524_),
    .X(_2545_));
 sky130_fd_sc_hd__clkbuf_1 _6217_ (.A(_2545_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _6218_ (.A0(net3),
    .A1(_0380_),
    .S(_2537_),
    .X(_2546_));
 sky130_fd_sc_hd__clkbuf_2 _6219_ (.A(_3095_),
    .X(_2547_));
 sky130_fd_sc_hd__and2_1 _6220_ (.A(_2546_),
    .B(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__clkbuf_1 _6221_ (.A(_2548_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _6222_ (.A0(net2),
    .A1(_0718_),
    .S(_2537_),
    .X(_2549_));
 sky130_fd_sc_hd__and2_1 _6223_ (.A(_2549_),
    .B(_2547_),
    .X(_2550_));
 sky130_fd_sc_hd__clkbuf_1 _6224_ (.A(_2550_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _6225_ (.A0(net16),
    .A1(_0385_),
    .S(_2537_),
    .X(_2551_));
 sky130_fd_sc_hd__and2_1 _6226_ (.A(_2551_),
    .B(_2547_),
    .X(_2552_));
 sky130_fd_sc_hd__clkbuf_1 _6227_ (.A(_2552_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _6228_ (.A0(net15),
    .A1(_0720_),
    .S(_2537_),
    .X(_2553_));
 sky130_fd_sc_hd__and2_1 _6229_ (.A(_2553_),
    .B(_2547_),
    .X(_2554_));
 sky130_fd_sc_hd__clkbuf_1 _6230_ (.A(_2554_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _6231_ (.A0(net14),
    .A1(_0868_),
    .S(_2537_),
    .X(_2555_));
 sky130_fd_sc_hd__and2_1 _6232_ (.A(_2555_),
    .B(_2547_),
    .X(_2556_));
 sky130_fd_sc_hd__clkbuf_1 _6233_ (.A(_2556_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _6234_ (.A0(net13),
    .A1(_0350_),
    .S(_2537_),
    .X(_2557_));
 sky130_fd_sc_hd__and2_1 _6235_ (.A(_2557_),
    .B(_2547_),
    .X(_2558_));
 sky130_fd_sc_hd__clkbuf_1 _6236_ (.A(_2558_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _6237_ (.A0(net12),
    .A1(_0337_),
    .S(_2536_),
    .X(_2559_));
 sky130_fd_sc_hd__and2_1 _6238_ (.A(_2559_),
    .B(_2547_),
    .X(_2560_));
 sky130_fd_sc_hd__clkbuf_1 _6239_ (.A(_2560_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _6240_ (.A0(net11),
    .A1(_0343_),
    .S(_2536_),
    .X(_2561_));
 sky130_fd_sc_hd__and2_1 _6241_ (.A(_2561_),
    .B(_2547_),
    .X(_2562_));
 sky130_fd_sc_hd__clkbuf_1 _6242_ (.A(_2562_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _6243_ (.A0(net10),
    .A1(_0408_),
    .S(_2536_),
    .X(_2563_));
 sky130_fd_sc_hd__and2_1 _6244_ (.A(_2563_),
    .B(_2547_),
    .X(_2564_));
 sky130_fd_sc_hd__clkbuf_1 _6245_ (.A(_2564_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _6246_ (.A0(net9),
    .A1(_0403_),
    .S(_2536_),
    .X(_2565_));
 sky130_fd_sc_hd__and2_1 _6247_ (.A(_2565_),
    .B(_2547_),
    .X(_2566_));
 sky130_fd_sc_hd__clkbuf_1 _6248_ (.A(_2566_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _6249_ (.A0(net8),
    .A1(_0392_),
    .S(_2536_),
    .X(_2567_));
 sky130_fd_sc_hd__buf_2 _6250_ (.A(_3095_),
    .X(_2568_));
 sky130_fd_sc_hd__and2_1 _6251_ (.A(_2567_),
    .B(_2568_),
    .X(_2569_));
 sky130_fd_sc_hd__clkbuf_1 _6252_ (.A(_2569_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _6253_ (.A0(net1),
    .A1(_0396_),
    .S(_2536_),
    .X(_2570_));
 sky130_fd_sc_hd__and2_1 _6254_ (.A(_2570_),
    .B(_2568_),
    .X(_2571_));
 sky130_fd_sc_hd__clkbuf_1 _6255_ (.A(_2571_),
    .X(_0200_));
 sky130_fd_sc_hd__or4b_1 _6256_ (.A(_3052_),
    .B(_3045_),
    .C(net41),
    .D_N(_3076_),
    .X(_2572_));
 sky130_fd_sc_hd__buf_2 _6257_ (.A(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_4 _6258_ (.A(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__mux2_1 _6259_ (.A0(net7),
    .A1(_0565_),
    .S(_2574_),
    .X(_2575_));
 sky130_fd_sc_hd__and2_1 _6260_ (.A(_2575_),
    .B(_2568_),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_1 _6261_ (.A(_2576_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _6262_ (.A0(net6),
    .A1(_0569_),
    .S(_2574_),
    .X(_2577_));
 sky130_fd_sc_hd__and2_1 _6263_ (.A(_2577_),
    .B(_2568_),
    .X(_2578_));
 sky130_fd_sc_hd__clkbuf_1 _6264_ (.A(_2578_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _6265_ (.A0(net5),
    .A1(_0580_),
    .S(_2574_),
    .X(_2579_));
 sky130_fd_sc_hd__and2_1 _6266_ (.A(_2579_),
    .B(_2568_),
    .X(_2580_));
 sky130_fd_sc_hd__clkbuf_1 _6267_ (.A(_2580_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _6268_ (.A0(net4),
    .A1(_0575_),
    .S(_2574_),
    .X(_2581_));
 sky130_fd_sc_hd__and2_1 _6269_ (.A(_2581_),
    .B(_2568_),
    .X(_2582_));
 sky130_fd_sc_hd__clkbuf_1 _6270_ (.A(_2582_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _6271_ (.A0(net3),
    .A1(_0590_),
    .S(_2574_),
    .X(_2583_));
 sky130_fd_sc_hd__and2_1 _6272_ (.A(_2583_),
    .B(_2568_),
    .X(_2584_));
 sky130_fd_sc_hd__clkbuf_1 _6273_ (.A(_2584_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _6274_ (.A0(net2),
    .A1(_0774_),
    .S(_2574_),
    .X(_2585_));
 sky130_fd_sc_hd__and2_1 _6275_ (.A(_2585_),
    .B(_2568_),
    .X(_2586_));
 sky130_fd_sc_hd__clkbuf_1 _6276_ (.A(_2586_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _6277_ (.A0(net16),
    .A1(_0595_),
    .S(_2574_),
    .X(_2587_));
 sky130_fd_sc_hd__and2_1 _6278_ (.A(_2587_),
    .B(_2568_),
    .X(_2588_));
 sky130_fd_sc_hd__clkbuf_1 _6279_ (.A(_2588_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _6280_ (.A0(net15),
    .A1(_0776_),
    .S(_2574_),
    .X(_2589_));
 sky130_fd_sc_hd__and2_1 _6281_ (.A(_2589_),
    .B(_2568_),
    .X(_2590_));
 sky130_fd_sc_hd__clkbuf_1 _6282_ (.A(_2590_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _6283_ (.A0(net14),
    .A1(_0561_),
    .S(_2574_),
    .X(_2591_));
 sky130_fd_sc_hd__buf_2 _6284_ (.A(net20),
    .X(_2592_));
 sky130_fd_sc_hd__and2_1 _6285_ (.A(_2591_),
    .B(_2592_),
    .X(_2593_));
 sky130_fd_sc_hd__clkbuf_1 _6286_ (.A(_2593_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _6287_ (.A0(net13),
    .A1(_0556_),
    .S(_2574_),
    .X(_2594_));
 sky130_fd_sc_hd__and2_1 _6288_ (.A(_2594_),
    .B(_2592_),
    .X(_2595_));
 sky130_fd_sc_hd__clkbuf_1 _6289_ (.A(_2595_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _6290_ (.A0(net12),
    .A1(_0542_),
    .S(_2573_),
    .X(_2596_));
 sky130_fd_sc_hd__and2_1 _6291_ (.A(_2596_),
    .B(_2592_),
    .X(_2597_));
 sky130_fd_sc_hd__clkbuf_1 _6292_ (.A(_2597_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _6293_ (.A0(net11),
    .A1(_0549_),
    .S(_2573_),
    .X(_2598_));
 sky130_fd_sc_hd__and2_1 _6294_ (.A(_2598_),
    .B(_2592_),
    .X(_2599_));
 sky130_fd_sc_hd__clkbuf_1 _6295_ (.A(_2599_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _6296_ (.A0(net10),
    .A1(_0602_),
    .S(_2573_),
    .X(_2600_));
 sky130_fd_sc_hd__and2_1 _6297_ (.A(_2600_),
    .B(_2592_),
    .X(_2601_));
 sky130_fd_sc_hd__clkbuf_1 _6298_ (.A(_2601_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _6299_ (.A0(net9),
    .A1(_0606_),
    .S(_2573_),
    .X(_2602_));
 sky130_fd_sc_hd__and2_1 _6300_ (.A(_2602_),
    .B(_2592_),
    .X(_2603_));
 sky130_fd_sc_hd__clkbuf_1 _6301_ (.A(_2603_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _6302_ (.A0(net8),
    .A1(_0781_),
    .S(_2573_),
    .X(_2604_));
 sky130_fd_sc_hd__and2_1 _6303_ (.A(_2604_),
    .B(_2592_),
    .X(_2605_));
 sky130_fd_sc_hd__clkbuf_1 _6304_ (.A(_2605_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _6305_ (.A0(net1),
    .A1(_0924_),
    .S(_2573_),
    .X(_2606_));
 sky130_fd_sc_hd__and2_1 _6306_ (.A(_2606_),
    .B(_2592_),
    .X(_2607_));
 sky130_fd_sc_hd__clkbuf_1 _6307_ (.A(_2607_),
    .X(_0184_));
 sky130_fd_sc_hd__or2_1 _6308_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .X(_2608_));
 sky130_fd_sc_hd__nand2_2 _6309_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2609_));
 sky130_fd_sc_hd__nand2_2 _6310_ (.A(_2608_),
    .B(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__o21ai_4 _6311_ (.A1(_3034_),
    .A2(_2610_),
    .B1(_2609_),
    .Y(_2611_));
 sky130_fd_sc_hd__or2_1 _6312_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .X(_2612_));
 sky130_fd_sc_hd__nand2_1 _6313_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2613_));
 sky130_fd_sc_hd__a21bo_2 _6314_ (.A1(_2611_),
    .A2(_2612_),
    .B1_N(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__o21ai_1 _6315_ (.A1(\egd_top.BitStream_buffer.pc_previous[3] ),
    .A2(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .B1(_2614_),
    .Y(_2615_));
 sky130_fd_sc_hd__nand2_1 _6316_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2616_));
 sky130_fd_sc_hd__nand2_2 _6317_ (.A(_2615_),
    .B(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__and3_2 _6318_ (.A(_2617_),
    .B(\egd_top.BitStream_buffer.pc_previous[4] ),
    .C(\egd_top.BitStream_buffer.pc_previous[5] ),
    .X(_2618_));
 sky130_fd_sc_hd__xor2_4 _6319_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_2618_),
    .X(\egd_top.BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(_3063_),
    .B(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2619_));
 sky130_fd_sc_hd__inv_2 _6321_ (.A(_2619_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21oi_1 _6322_ (.A1(_2617_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[5] ),
    .Y(_2620_));
 sky130_fd_sc_hd__nor2_2 _6323_ (.A(_2620_),
    .B(_2618_),
    .Y(\egd_top.BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__nand2_1 _6324_ (.A(_3063_),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_2621_));
 sky130_fd_sc_hd__inv_2 _6325_ (.A(_2621_),
    .Y(_0182_));
 sky130_fd_sc_hd__xor2_4 _6326_ (.A(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B(_2617_),
    .X(\egd_top.BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__nand2_1 _6327_ (.A(_3063_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_2622_));
 sky130_fd_sc_hd__inv_2 _6328_ (.A(_2622_),
    .Y(_0181_));
 sky130_fd_sc_hd__nor2_1 _6329_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2623_));
 sky130_fd_sc_hd__and2b_2 _6330_ (.A_N(_2623_),
    .B(_2616_),
    .X(_2624_));
 sky130_fd_sc_hd__xor2_4 _6331_ (.A(_2624_),
    .B(_2614_),
    .X(\egd_top.BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__nand2_1 _6332_ (.A(_3063_),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2625_));
 sky130_fd_sc_hd__inv_2 _6333_ (.A(_2625_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_2 _6334_ (.A(_2612_),
    .B(_2613_),
    .Y(_2626_));
 sky130_fd_sc_hd__xnor2_4 _6335_ (.A(_2626_),
    .B(_2611_),
    .Y(\egd_top.BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__nand2_1 _6336_ (.A(_3063_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_2627_));
 sky130_fd_sc_hd__inv_2 _6337_ (.A(_2627_),
    .Y(_0179_));
 sky130_fd_sc_hd__xor2_4 _6338_ (.A(_3034_),
    .B(_2610_),
    .X(\egd_top.BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__nand2_1 _6339_ (.A(_3063_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2628_));
 sky130_fd_sc_hd__inv_2 _6340_ (.A(_2628_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_1 _6341_ (.A(_3036_),
    .B(_3063_),
    .Y(_2629_));
 sky130_fd_sc_hd__inv_2 _6342_ (.A(_2629_),
    .Y(_0177_));
 sky130_fd_sc_hd__or4b_1 _6343_ (.A(_3052_),
    .B(net39),
    .C(_3046_),
    .D_N(_3076_),
    .X(_2630_));
 sky130_fd_sc_hd__buf_2 _6344_ (.A(net40),
    .X(_2631_));
 sky130_fd_sc_hd__clkbuf_4 _6345_ (.A(_2631_),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_1 _6346_ (.A0(net7),
    .A1(_0725_),
    .S(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__and2_1 _6347_ (.A(_2633_),
    .B(_2592_),
    .X(_2634_));
 sky130_fd_sc_hd__clkbuf_1 _6348_ (.A(_2634_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _6349_ (.A0(net6),
    .A1(_0872_),
    .S(_2632_),
    .X(_2635_));
 sky130_fd_sc_hd__and2_1 _6350_ (.A(_2635_),
    .B(_2592_),
    .X(_2636_));
 sky130_fd_sc_hd__clkbuf_1 _6351_ (.A(_2636_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _6352_ (.A0(net5),
    .A1(_0749_),
    .S(_2632_),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_2 _6353_ (.A(net20),
    .X(_2638_));
 sky130_fd_sc_hd__and2_1 _6354_ (.A(_2637_),
    .B(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _6355_ (.A(_2639_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _6356_ (.A0(net4),
    .A1(_0500_),
    .S(_2632_),
    .X(_2640_));
 sky130_fd_sc_hd__and2_1 _6357_ (.A(_2640_),
    .B(_2638_),
    .X(_2641_));
 sky130_fd_sc_hd__clkbuf_1 _6358_ (.A(_2641_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _6359_ (.A0(net3),
    .A1(_0751_),
    .S(_2632_),
    .X(_2642_));
 sky130_fd_sc_hd__and2_1 _6360_ (.A(_2642_),
    .B(_2638_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _6361_ (.A(_2643_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _6362_ (.A0(net2),
    .A1(_0897_),
    .S(_2632_),
    .X(_2644_));
 sky130_fd_sc_hd__and2_1 _6363_ (.A(_2644_),
    .B(_2638_),
    .X(_2645_));
 sky130_fd_sc_hd__clkbuf_1 _6364_ (.A(_2645_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _6365_ (.A0(net16),
    .A1(_1032_),
    .S(_2632_),
    .X(_2646_));
 sky130_fd_sc_hd__and2_1 _6366_ (.A(_2646_),
    .B(_2638_),
    .X(_2647_));
 sky130_fd_sc_hd__clkbuf_1 _6367_ (.A(_2647_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _6368_ (.A0(net15),
    .A1(_0522_),
    .S(_2632_),
    .X(_2648_));
 sky130_fd_sc_hd__and2_1 _6369_ (.A(_2648_),
    .B(_2638_),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_1 _6370_ (.A(_2649_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _6371_ (.A0(net14),
    .A1(_0758_),
    .S(_2632_),
    .X(_2650_));
 sky130_fd_sc_hd__and2_1 _6372_ (.A(_2650_),
    .B(_2638_),
    .X(_2651_));
 sky130_fd_sc_hd__clkbuf_1 _6373_ (.A(_2651_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _6374_ (.A0(net13),
    .A1(_0904_),
    .S(_2632_),
    .X(_2652_));
 sky130_fd_sc_hd__and2_1 _6375_ (.A(_2652_),
    .B(_2638_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_1 _6376_ (.A(_2653_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _6377_ (.A0(net12),
    .A1(_0474_),
    .S(_2631_),
    .X(_2654_));
 sky130_fd_sc_hd__and2_1 _6378_ (.A(_2654_),
    .B(_2638_),
    .X(_2655_));
 sky130_fd_sc_hd__clkbuf_1 _6379_ (.A(_2655_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _6380_ (.A0(net11),
    .A1(_0481_),
    .S(_2631_),
    .X(_2656_));
 sky130_fd_sc_hd__and2_1 _6381_ (.A(_2656_),
    .B(_2638_),
    .X(_2657_));
 sky130_fd_sc_hd__clkbuf_1 _6382_ (.A(_2657_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _6383_ (.A0(net10),
    .A1(_0745_),
    .S(_2631_),
    .X(_2658_));
 sky130_fd_sc_hd__and2_1 _6384_ (.A(_2658_),
    .B(_3008_),
    .X(_2659_));
 sky130_fd_sc_hd__clkbuf_1 _6385_ (.A(_2659_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _6386_ (.A0(net9),
    .A1(_0892_),
    .S(_2631_),
    .X(_2660_));
 sky130_fd_sc_hd__and2_1 _6387_ (.A(_2660_),
    .B(_3008_),
    .X(_2661_));
 sky130_fd_sc_hd__clkbuf_1 _6388_ (.A(_2661_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _6389_ (.A0(net8),
    .A1(_0525_),
    .S(_2631_),
    .X(_2662_));
 sky130_fd_sc_hd__and2_1 _6390_ (.A(_2662_),
    .B(_3008_),
    .X(_2663_));
 sky130_fd_sc_hd__clkbuf_1 _6391_ (.A(_2663_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _6392_ (.A0(net1),
    .A1(_0529_),
    .S(_2631_),
    .X(_2664_));
 sky130_fd_sc_hd__and2_1 _6393_ (.A(_2664_),
    .B(_3008_),
    .X(_2665_));
 sky130_fd_sc_hd__clkbuf_1 _6394_ (.A(_2665_),
    .X(_0161_));
 sky130_fd_sc_hd__inv_2 _6395_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2666_));
 sky130_fd_sc_hd__nand2_1 _6396_ (.A(_2666_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2667_));
 sky130_fd_sc_hd__inv_2 _6397_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2668_));
 sky130_fd_sc_hd__nand2_1 _6398_ (.A(_2667_),
    .B(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__inv_2 _6399_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2670_));
 sky130_fd_sc_hd__nand2_1 _6400_ (.A(_2669_),
    .B(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__inv_2 _6401_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2672_));
 sky130_fd_sc_hd__nand2_1 _6402_ (.A(_2671_),
    .B(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__inv_2 _6403_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2674_));
 sky130_fd_sc_hd__nand2_1 _6404_ (.A(_2673_),
    .B(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__inv_2 _6405_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2676_));
 sky130_fd_sc_hd__nand2_1 _6406_ (.A(_2675_),
    .B(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__inv_2 _6407_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_2678_));
 sky130_fd_sc_hd__nand2_1 _6408_ (.A(_2677_),
    .B(_2678_),
    .Y(_2679_));
 sky130_fd_sc_hd__inv_2 _6409_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2680_));
 sky130_fd_sc_hd__nand2_1 _6410_ (.A(_2679_),
    .B(_2680_),
    .Y(_2681_));
 sky130_fd_sc_hd__inv_2 _6411_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2682_));
 sky130_fd_sc_hd__inv_4 _6412_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2683_));
 sky130_fd_sc_hd__nand2_1 _6413_ (.A(_2682_),
    .B(_2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__nor2_1 _6414_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(_2684_),
    .Y(_2685_));
 sky130_fd_sc_hd__inv_2 _6415_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_2686_));
 sky130_fd_sc_hd__nand2_1 _6416_ (.A(_2685_),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__inv_2 _6417_ (.A(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__nand2_1 _6418_ (.A(_2681_),
    .B(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__a21oi_1 _6419_ (.A1(_2682_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2690_));
 sky130_fd_sc_hd__nand2_1 _6420_ (.A(_2689_),
    .B(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__nor2_1 _6421_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2692_));
 sky130_fd_sc_hd__nand2_1 _6422_ (.A(_2691_),
    .B(_2692_),
    .Y(_2693_));
 sky130_fd_sc_hd__nor2_1 _6423_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_2694_));
 sky130_fd_sc_hd__nand2_2 _6424_ (.A(_2693_),
    .B(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__and3_1 _6425_ (.A(_2688_),
    .B(_2680_),
    .C(_2678_),
    .X(_2696_));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(_2692_),
    .B(_3070_),
    .Y(_2697_));
 sky130_fd_sc_hd__inv_2 _6427_ (.A(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__and2_1 _6428_ (.A(_2696_),
    .B(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__nor2_1 _6429_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2700_));
 sky130_fd_sc_hd__inv_2 _6430_ (.A(_2700_),
    .Y(_2701_));
 sky130_fd_sc_hd__nor2_1 _6431_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2701_),
    .Y(_2702_));
 sky130_fd_sc_hd__nand2_1 _6432_ (.A(_2702_),
    .B(_2670_),
    .Y(_2703_));
 sky130_fd_sc_hd__nor2_1 _6433_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2704_));
 sky130_fd_sc_hd__nand2_1 _6434_ (.A(_2698_),
    .B(_2704_),
    .Y(_2705_));
 sky130_fd_sc_hd__a21o_1 _6435_ (.A1(_2696_),
    .A2(_2703_),
    .B1(_2705_),
    .X(_2706_));
 sky130_fd_sc_hd__nor2_1 _6436_ (.A(_2699_),
    .B(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__o21a_1 _6437_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_2670_),
    .X(_2708_));
 sky130_fd_sc_hd__a211o_1 _6438_ (.A1(_2708_),
    .A2(_2672_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .C1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .X(_2709_));
 sky130_fd_sc_hd__a21o_1 _6439_ (.A1(_2687_),
    .A2(_2704_),
    .B1(_2697_),
    .X(_2710_));
 sky130_fd_sc_hd__a21oi_2 _6440_ (.A1(_2709_),
    .A2(_2696_),
    .B1(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__inv_2 _6441_ (.A(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__nand3b_2 _6442_ (.A_N(_2695_),
    .B(_2707_),
    .C(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hd__nor2_1 _6443_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .B(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(_2711_),
    .B(_2705_),
    .Y(_2715_));
 sky130_fd_sc_hd__a21oi_1 _6445_ (.A1(_2693_),
    .A2(_2694_),
    .B1(_2715_),
    .Y(_2716_));
 sky130_fd_sc_hd__inv_2 _6446_ (.A(_2707_),
    .Y(_2717_));
 sky130_fd_sc_hd__buf_6 _6447_ (.A(_2717_),
    .X(_2718_));
 sky130_fd_sc_hd__nor2_1 _6448_ (.A(_2711_),
    .B(_2718_),
    .Y(_2719_));
 sky130_fd_sc_hd__nand2_2 _6449_ (.A(_2719_),
    .B(_2695_),
    .Y(_2720_));
 sky130_fd_sc_hd__o2bb2ai_1 _6450_ (.A1_N(_2683_),
    .A2_N(_2716_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B2(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__nor2_1 _6451_ (.A(_2714_),
    .B(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__nand3_1 _6452_ (.A(_2693_),
    .B(_2711_),
    .C(_2694_),
    .Y(_2723_));
 sky130_fd_sc_hd__buf_4 _6453_ (.A(_2723_),
    .X(_2724_));
 sky130_fd_sc_hd__o21ai_1 _6454_ (.A1(_2718_),
    .A2(_2724_),
    .B1(_2668_),
    .Y(_2725_));
 sky130_fd_sc_hd__nor2_1 _6455_ (.A(_2717_),
    .B(_2723_),
    .Y(_2726_));
 sky130_fd_sc_hd__buf_6 _6456_ (.A(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__inv_2 _6457_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2728_));
 sky130_fd_sc_hd__nand2_1 _6458_ (.A(_2727_),
    .B(_2728_),
    .Y(_2729_));
 sky130_fd_sc_hd__nand2_1 _6459_ (.A(_2725_),
    .B(_2729_),
    .Y(_2730_));
 sky130_fd_sc_hd__nor2_2 _6460_ (.A(_2712_),
    .B(_2718_),
    .Y(_2731_));
 sky130_fd_sc_hd__nand2_1 _6461_ (.A(_2730_),
    .B(_2731_),
    .Y(_2732_));
 sky130_fd_sc_hd__inv_2 _6462_ (.A(_2705_),
    .Y(_2733_));
 sky130_fd_sc_hd__nor2_1 _6463_ (.A(_2733_),
    .B(_2724_),
    .Y(_2734_));
 sky130_fd_sc_hd__nor3_1 _6464_ (.A(_2733_),
    .B(_2711_),
    .C(_2695_),
    .Y(_2735_));
 sky130_fd_sc_hd__inv_2 _6465_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2736_));
 sky130_fd_sc_hd__a22oi_2 _6466_ (.A1(_2734_),
    .A2(_2680_),
    .B1(_2735_),
    .B2(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__nand3_2 _6467_ (.A(_2722_),
    .B(_2732_),
    .C(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__nand2_4 _6468_ (.A(_2738_),
    .B(_3032_),
    .Y(_2739_));
 sky130_fd_sc_hd__inv_2 _6469_ (.A(_3032_),
    .Y(_2740_));
 sky130_fd_sc_hd__a311o_1 _6470_ (.A1(_2695_),
    .A2(_2712_),
    .A3(_2706_),
    .B1(_2740_),
    .C1(_2699_),
    .X(_2741_));
 sky130_fd_sc_hd__nand2_1 _6471_ (.A(net18),
    .B(net17),
    .Y(_2742_));
 sky130_fd_sc_hd__inv_2 _6472_ (.A(_2742_),
    .Y(_2743_));
 sky130_fd_sc_hd__and3b_1 _6473_ (.A_N(net23),
    .B(_2743_),
    .C(net22),
    .X(_2744_));
 sky130_fd_sc_hd__inv_2 _6474_ (.A(\egd_top.exp_golomb_decoding.te_range[2] ),
    .Y(_2745_));
 sky130_fd_sc_hd__and2_2 _6475_ (.A(_2744_),
    .B(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__inv_4 _6476_ (.A(_2739_),
    .Y(_2747_));
 sky130_fd_sc_hd__nor2_1 _6477_ (.A(_2746_),
    .B(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__a211o_1 _6478_ (.A1(_2741_),
    .A2(_2746_),
    .B1(_2742_),
    .C1(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__nor2_2 _6479_ (.A(net17),
    .B(_3030_),
    .Y(_2750_));
 sky130_fd_sc_hd__inv_2 _6480_ (.A(_2750_),
    .Y(_2751_));
 sky130_fd_sc_hd__xnor2_1 _6481_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2752_));
 sky130_fd_sc_hd__nand2_1 _6482_ (.A(_2735_),
    .B(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__nor2_1 _6483_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2754_));
 sky130_fd_sc_hd__inv_2 _6484_ (.A(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__nand2_1 _6485_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2756_));
 sky130_fd_sc_hd__nand2_1 _6486_ (.A(_2755_),
    .B(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__nand2_1 _6487_ (.A(_2734_),
    .B(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__nand2_1 _6488_ (.A(_2753_),
    .B(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__inv_2 _6489_ (.A(_2713_),
    .Y(_2760_));
 sky130_fd_sc_hd__nand2_1 _6490_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2761_));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(_2701_),
    .B(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__nand2_1 _6492_ (.A(_2760_),
    .B(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__inv_2 _6493_ (.A(_2720_),
    .Y(_2764_));
 sky130_fd_sc_hd__nor2_1 _6494_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2765_));
 sky130_fd_sc_hd__inv_2 _6495_ (.A(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__nand2_1 _6496_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2767_));
 sky130_fd_sc_hd__nand2_1 _6497_ (.A(_2766_),
    .B(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__nand2_1 _6498_ (.A(_2764_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__xnor2_1 _6499_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2770_));
 sky130_fd_sc_hd__nand2_1 _6500_ (.A(_2716_),
    .B(_2770_),
    .Y(_2771_));
 sky130_fd_sc_hd__nand3_1 _6501_ (.A(_2763_),
    .B(_2769_),
    .C(_2771_),
    .Y(_2772_));
 sky130_fd_sc_hd__nor2_1 _6502_ (.A(_2759_),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__nand2_1 _6503_ (.A(_2726_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2774_));
 sky130_fd_sc_hd__o21ai_1 _6504_ (.A1(_2670_),
    .A2(_2727_),
    .B1(_2774_),
    .Y(_2775_));
 sky130_fd_sc_hd__nand2_1 _6505_ (.A(_2775_),
    .B(_2730_),
    .Y(_2776_));
 sky130_fd_sc_hd__o21ai_1 _6506_ (.A1(_2718_),
    .A2(_2724_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2777_));
 sky130_fd_sc_hd__nand2_1 _6507_ (.A(_2726_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2778_));
 sky130_fd_sc_hd__nand2_1 _6508_ (.A(_2777_),
    .B(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__o21ai_1 _6509_ (.A1(_2718_),
    .A2(_2724_),
    .B1(_2670_),
    .Y(_2780_));
 sky130_fd_sc_hd__inv_2 _6510_ (.A(_2724_),
    .Y(_2781_));
 sky130_fd_sc_hd__nand3_1 _6511_ (.A(_2781_),
    .B(_2666_),
    .C(_2707_),
    .Y(_2782_));
 sky130_fd_sc_hd__nand2_1 _6512_ (.A(_2780_),
    .B(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__nand2_1 _6513_ (.A(_2779_),
    .B(_2783_),
    .Y(_2784_));
 sky130_fd_sc_hd__nand3_1 _6514_ (.A(_2776_),
    .B(_2784_),
    .C(_2731_),
    .Y(_2785_));
 sky130_fd_sc_hd__nand2_1 _6515_ (.A(_2773_),
    .B(_2785_),
    .Y(_2786_));
 sky130_fd_sc_hd__buf_4 _6516_ (.A(_3032_),
    .X(_2787_));
 sky130_fd_sc_hd__nand2_1 _6517_ (.A(_2786_),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__inv_2 _6518_ (.A(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__nor2_1 _6519_ (.A(_2747_),
    .B(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__nand3_1 _6520_ (.A(_2786_),
    .B(_2738_),
    .C(_2787_),
    .Y(_2791_));
 sky130_fd_sc_hd__or3b_1 _6521_ (.A(_2751_),
    .B(_2790_),
    .C_N(_2791_),
    .X(_2792_));
 sky130_fd_sc_hd__o311ai_4 _6522_ (.A1(net18),
    .A2(_3031_),
    .A3(_2739_),
    .B1(_2749_),
    .C1(_2792_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_1 _6523_ (.A(_2730_),
    .B(_2783_),
    .Y(_2793_));
 sky130_fd_sc_hd__o21ai_1 _6524_ (.A1(_2718_),
    .A2(_2724_),
    .B1(_2672_),
    .Y(_2794_));
 sky130_fd_sc_hd__nand2_1 _6525_ (.A(_2727_),
    .B(_2668_),
    .Y(_2795_));
 sky130_fd_sc_hd__nand2_1 _6526_ (.A(_2794_),
    .B(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__nand2_1 _6527_ (.A(_2793_),
    .B(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__o21ai_1 _6528_ (.A1(_2718_),
    .A2(_2724_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2798_));
 sky130_fd_sc_hd__nand2_1 _6529_ (.A(_2727_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2799_));
 sky130_fd_sc_hd__nand2_1 _6530_ (.A(_2798_),
    .B(_2799_),
    .Y(_2800_));
 sky130_fd_sc_hd__nand3_1 _6531_ (.A(_2730_),
    .B(_2800_),
    .C(_2783_),
    .Y(_2801_));
 sky130_fd_sc_hd__nand3_1 _6532_ (.A(_2797_),
    .B(_2801_),
    .C(_2731_),
    .Y(_2802_));
 sky130_fd_sc_hd__nor2_1 _6533_ (.A(_2680_),
    .B(_2765_),
    .Y(_2803_));
 sky130_fd_sc_hd__nor2_1 _6534_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2766_),
    .Y(_2804_));
 sky130_fd_sc_hd__nor2_1 _6535_ (.A(_2803_),
    .B(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__and2_1 _6536_ (.A(_2684_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .X(_2806_));
 sky130_fd_sc_hd__o21ai_1 _6537_ (.A1(_2685_),
    .A2(_2806_),
    .B1(_2716_),
    .Y(_2807_));
 sky130_fd_sc_hd__o21ai_1 _6538_ (.A1(_2805_),
    .A2(_2720_),
    .B1(_2807_),
    .Y(_2808_));
 sky130_fd_sc_hd__nor2_1 _6539_ (.A(_2676_),
    .B(_2700_),
    .Y(_2809_));
 sky130_fd_sc_hd__nor2_1 _6540_ (.A(_2809_),
    .B(_2702_),
    .Y(_2810_));
 sky130_fd_sc_hd__nor2_1 _6541_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2755_),
    .Y(_2811_));
 sky130_fd_sc_hd__nor2_1 _6542_ (.A(_2683_),
    .B(_2754_),
    .Y(_2812_));
 sky130_fd_sc_hd__o21ai_1 _6543_ (.A1(_2811_),
    .A2(_2812_),
    .B1(_2734_),
    .Y(_2813_));
 sky130_fd_sc_hd__o21ai_1 _6544_ (.A1(_2810_),
    .A2(_2713_),
    .B1(_2813_),
    .Y(_2814_));
 sky130_fd_sc_hd__nor2_1 _6545_ (.A(_2808_),
    .B(_2814_),
    .Y(_2815_));
 sky130_fd_sc_hd__nand2_1 _6546_ (.A(_2802_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__nand2_2 _6547_ (.A(_2816_),
    .B(_2787_),
    .Y(_2817_));
 sky130_fd_sc_hd__or2_1 _6548_ (.A(_2788_),
    .B(_2817_),
    .X(_2818_));
 sky130_fd_sc_hd__nand2_1 _6549_ (.A(_2817_),
    .B(_2788_),
    .Y(_2819_));
 sky130_fd_sc_hd__a31o_1 _6550_ (.A1(_2744_),
    .A2(net18),
    .A3(_2745_),
    .B1(_3031_),
    .X(_2820_));
 sky130_fd_sc_hd__inv_2 _6551_ (.A(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__a32o_1 _6552_ (.A1(_2818_),
    .A2(_2819_),
    .A3(_2750_),
    .B1(_2789_),
    .B2(_2821_),
    .X(net23));
 sky130_fd_sc_hd__o21ai_1 _6553_ (.A1(_2788_),
    .A2(_2817_),
    .B1(_2747_),
    .Y(_2822_));
 sky130_fd_sc_hd__nand2_1 _6554_ (.A(_2822_),
    .B(_2819_),
    .Y(_2823_));
 sky130_fd_sc_hd__nor2_1 _6555_ (.A(_2779_),
    .B(_2775_),
    .Y(_2824_));
 sky130_fd_sc_hd__o21ai_1 _6556_ (.A1(_2718_),
    .A2(_2724_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2825_));
 sky130_fd_sc_hd__nand2_1 _6557_ (.A(_2726_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2826_));
 sky130_fd_sc_hd__nand2_1 _6558_ (.A(_2825_),
    .B(_2826_),
    .Y(_2827_));
 sky130_fd_sc_hd__nand3_1 _6559_ (.A(_2824_),
    .B(_2827_),
    .C(_2796_),
    .Y(_2828_));
 sky130_fd_sc_hd__nand3_1 _6560_ (.A(_2730_),
    .B(_2796_),
    .C(_2783_),
    .Y(_2829_));
 sky130_fd_sc_hd__nand2_1 _6561_ (.A(_2727_),
    .B(_2670_),
    .Y(_2830_));
 sky130_fd_sc_hd__o21ai_1 _6562_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .A2(_2727_),
    .B1(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_1 _6563_ (.A(_2829_),
    .B(_2831_),
    .Y(_2832_));
 sky130_fd_sc_hd__nand3_1 _6564_ (.A(_2828_),
    .B(_2731_),
    .C(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__nor2_1 _6565_ (.A(_2701_),
    .B(_2766_),
    .Y(_2834_));
 sky130_fd_sc_hd__nor2_1 _6566_ (.A(_2678_),
    .B(_2702_),
    .Y(_2835_));
 sky130_fd_sc_hd__o21ai_1 _6567_ (.A1(_2834_),
    .A2(_2835_),
    .B1(_2760_),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_1 _6568_ (.A(_2684_),
    .B(_2755_),
    .Y(_2837_));
 sky130_fd_sc_hd__nor2_1 _6569_ (.A(_2682_),
    .B(_2811_),
    .Y(_2838_));
 sky130_fd_sc_hd__o21ai_1 _6570_ (.A1(_2837_),
    .A2(_2838_),
    .B1(_2734_),
    .Y(_2839_));
 sky130_fd_sc_hd__mux2_1 _6571_ (.A0(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .A1(_2757_),
    .S(_2765_),
    .X(_2840_));
 sky130_fd_sc_hd__nand2_1 _6572_ (.A(_2764_),
    .B(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__and3_1 _6573_ (.A(_2836_),
    .B(_2839_),
    .C(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__a21oi_1 _6574_ (.A1(_2833_),
    .A2(_2842_),
    .B1(_2740_),
    .Y(_2843_));
 sky130_fd_sc_hd__nand2_1 _6575_ (.A(_2823_),
    .B(_2843_),
    .Y(_2844_));
 sky130_fd_sc_hd__nand2_1 _6576_ (.A(_2833_),
    .B(_2842_),
    .Y(_2845_));
 sky130_fd_sc_hd__nand2_1 _6577_ (.A(_2845_),
    .B(_2787_),
    .Y(_2846_));
 sky130_fd_sc_hd__nand3_1 _6578_ (.A(_2822_),
    .B(_2819_),
    .C(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__nand2_1 _6579_ (.A(_2844_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__nand2_1 _6580_ (.A(_2848_),
    .B(_2750_),
    .Y(_2849_));
 sky130_fd_sc_hd__or2_1 _6581_ (.A(_2820_),
    .B(_2817_),
    .X(_2850_));
 sky130_fd_sc_hd__nand2_1 _6582_ (.A(net22),
    .B(net23),
    .Y(_2851_));
 sky130_fd_sc_hd__a21oi_1 _6583_ (.A1(_2849_),
    .A2(_2850_),
    .B1(_2851_),
    .Y(_2852_));
 sky130_fd_sc_hd__nand3_1 _6584_ (.A(_2849_),
    .B(_2851_),
    .C(_2850_),
    .Y(_2853_));
 sky130_fd_sc_hd__nand2_1 _6585_ (.A(_2853_),
    .B(_2743_),
    .Y(_2854_));
 sky130_fd_sc_hd__nor2_1 _6586_ (.A(_2852_),
    .B(_2854_),
    .Y(\egd_top.exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__or3_1 _6587_ (.A(_2740_),
    .B(_2746_),
    .C(_2695_),
    .X(_2855_));
 sky130_fd_sc_hd__inv_2 _6588_ (.A(_2855_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__or3_1 _6589_ (.A(_2740_),
    .B(_2746_),
    .C(_2712_),
    .X(_2856_));
 sky130_fd_sc_hd__inv_2 _6590_ (.A(_2856_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__or3_1 _6591_ (.A(_2740_),
    .B(_2746_),
    .C(_2706_),
    .X(_2857_));
 sky130_fd_sc_hd__inv_2 _6592_ (.A(_2857_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__nand2_1 _6593_ (.A(_2849_),
    .B(_2850_),
    .Y(net24));
 sky130_fd_sc_hd__nor2_1 _6594_ (.A(_2819_),
    .B(_2843_),
    .Y(_2858_));
 sky130_fd_sc_hd__nand2_1 _6595_ (.A(_2858_),
    .B(_2739_),
    .Y(_2859_));
 sky130_fd_sc_hd__nor2_1 _6596_ (.A(_2817_),
    .B(_2791_),
    .Y(_2860_));
 sky130_fd_sc_hd__nand2_1 _6597_ (.A(_2843_),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__nand2_1 _6598_ (.A(_2861_),
    .B(_2747_),
    .Y(_2862_));
 sky130_fd_sc_hd__nand2_1 _6599_ (.A(_2831_),
    .B(_2796_),
    .Y(_2863_));
 sky130_fd_sc_hd__o21ai_1 _6600_ (.A1(_2718_),
    .A2(_2724_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2864_));
 sky130_fd_sc_hd__nand2_1 _6601_ (.A(_2727_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2865_));
 sky130_fd_sc_hd__nand2_1 _6602_ (.A(_2864_),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__inv_2 _6603_ (.A(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__o21ai_1 _6604_ (.A1(_2793_),
    .A2(_2863_),
    .B1(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__nor2_1 _6605_ (.A(_2827_),
    .B(_2800_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand3_1 _6606_ (.A(_2824_),
    .B(_2869_),
    .C(_2866_),
    .Y(_2870_));
 sky130_fd_sc_hd__nand3_1 _6607_ (.A(_2868_),
    .B(_2870_),
    .C(_2731_),
    .Y(_2871_));
 sky130_fd_sc_hd__nand2_1 _6608_ (.A(_2765_),
    .B(_2754_),
    .Y(_2872_));
 sky130_fd_sc_hd__and2_1 _6609_ (.A(_2872_),
    .B(_2683_),
    .X(_2873_));
 sky130_fd_sc_hd__nor2_1 _6610_ (.A(_2683_),
    .B(_2872_),
    .Y(_2874_));
 sky130_fd_sc_hd__inv_2 _6611_ (.A(_2834_),
    .Y(_2875_));
 sky130_fd_sc_hd__nor2_1 _6612_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__nor2_1 _6613_ (.A(_2680_),
    .B(_2834_),
    .Y(_2877_));
 sky130_fd_sc_hd__o21ai_1 _6614_ (.A1(_2876_),
    .A2(_2877_),
    .B1(_2760_),
    .Y(_2878_));
 sky130_fd_sc_hd__o31a_1 _6615_ (.A1(_2873_),
    .A2(_2720_),
    .A3(_2874_),
    .B1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a21oi_1 _6616_ (.A1(_2871_),
    .A2(_2879_),
    .B1(_2740_),
    .Y(_2880_));
 sky130_fd_sc_hd__a21oi_1 _6617_ (.A1(_2859_),
    .A2(_2862_),
    .B1(_2880_),
    .Y(_2881_));
 sky130_fd_sc_hd__nand3_1 _6618_ (.A(_2859_),
    .B(_2862_),
    .C(_2880_),
    .Y(_2882_));
 sky130_fd_sc_hd__nand2_1 _6619_ (.A(_2882_),
    .B(_2750_),
    .Y(_2883_));
 sky130_fd_sc_hd__o2bb2ai_2 _6620_ (.A1_N(_2845_),
    .A2_N(_2821_),
    .B1(_2881_),
    .B2(_2883_),
    .Y(net25));
 sky130_fd_sc_hd__nand2_1 _6621_ (.A(_2871_),
    .B(_2879_),
    .Y(_2884_));
 sky130_fd_sc_hd__nand2_1 _6622_ (.A(_2884_),
    .B(_2787_),
    .Y(_2885_));
 sky130_fd_sc_hd__o21ai_1 _6623_ (.A1(_2885_),
    .A2(_2861_),
    .B1(_2747_),
    .Y(_2886_));
 sky130_fd_sc_hd__o21bai_1 _6624_ (.A1(_2786_),
    .A2(_2816_),
    .B1_N(_2740_),
    .Y(_2887_));
 sky130_fd_sc_hd__nand2_1 _6625_ (.A(_2887_),
    .B(_2846_),
    .Y(_2888_));
 sky130_fd_sc_hd__nor2_1 _6626_ (.A(_2880_),
    .B(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__nand2_1 _6627_ (.A(_2889_),
    .B(_2739_),
    .Y(_2890_));
 sky130_fd_sc_hd__nand2_1 _6628_ (.A(_2886_),
    .B(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__nand3_1 _6629_ (.A(_2824_),
    .B(_2869_),
    .C(_2867_),
    .Y(_2892_));
 sky130_fd_sc_hd__o21ai_1 _6630_ (.A1(_2718_),
    .A2(_2724_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_2893_));
 sky130_fd_sc_hd__nand2_1 _6631_ (.A(_2727_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2894_));
 sky130_fd_sc_hd__nand2_1 _6632_ (.A(_2893_),
    .B(_2894_),
    .Y(_2895_));
 sky130_fd_sc_hd__inv_2 _6633_ (.A(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__nand2_1 _6634_ (.A(_2892_),
    .B(_2896_),
    .Y(_2897_));
 sky130_fd_sc_hd__nor2_1 _6635_ (.A(_2793_),
    .B(_2863_),
    .Y(_2898_));
 sky130_fd_sc_hd__nand3_1 _6636_ (.A(_2898_),
    .B(_2895_),
    .C(_2867_),
    .Y(_2899_));
 sky130_fd_sc_hd__nand3_1 _6637_ (.A(_2897_),
    .B(_2899_),
    .C(_2731_),
    .Y(_2900_));
 sky130_fd_sc_hd__nor2_1 _6638_ (.A(_2757_),
    .B(_2875_),
    .Y(_2901_));
 sky130_fd_sc_hd__a211o_1 _6639_ (.A1(_2686_),
    .A2(_2875_),
    .B1(_2901_),
    .C1(_2713_),
    .X(_2902_));
 sky130_fd_sc_hd__nand2_1 _6640_ (.A(_2900_),
    .B(_2902_),
    .Y(_2903_));
 sky130_fd_sc_hd__nand2_1 _6641_ (.A(_2903_),
    .B(_2787_),
    .Y(_2904_));
 sky130_fd_sc_hd__nand2_1 _6642_ (.A(_2891_),
    .B(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__nand3b_1 _6643_ (.A_N(_2904_),
    .B(_2886_),
    .C(_2890_),
    .Y(_2906_));
 sky130_fd_sc_hd__nand3_1 _6644_ (.A(_2905_),
    .B(_2906_),
    .C(_2750_),
    .Y(_2907_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(_2884_),
    .B(_2821_),
    .Y(_2908_));
 sky130_fd_sc_hd__nand2_1 _6646_ (.A(_2907_),
    .B(_2908_),
    .Y(net26));
 sky130_fd_sc_hd__nand3_1 _6647_ (.A(_2903_),
    .B(_2787_),
    .C(_2884_),
    .Y(_2909_));
 sky130_fd_sc_hd__inv_2 _6648_ (.A(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__nor3_1 _6649_ (.A(_2817_),
    .B(_2791_),
    .C(_2846_),
    .Y(_2911_));
 sky130_fd_sc_hd__nand2_1 _6650_ (.A(_2910_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__inv_2 _6651_ (.A(_2731_),
    .Y(_2913_));
 sky130_fd_sc_hd__nor2_1 _6652_ (.A(_2895_),
    .B(_2866_),
    .Y(_2914_));
 sky130_fd_sc_hd__nand3_1 _6653_ (.A(_2824_),
    .B(_2914_),
    .C(_2869_),
    .Y(_2915_));
 sky130_fd_sc_hd__a21o_1 _6654_ (.A1(_2727_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .X(_2916_));
 sky130_fd_sc_hd__inv_2 _6655_ (.A(_2916_),
    .Y(_2917_));
 sky130_fd_sc_hd__nand2_1 _6656_ (.A(_2915_),
    .B(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__nand3_1 _6657_ (.A(_2898_),
    .B(_2914_),
    .C(_2916_),
    .Y(_2919_));
 sky130_fd_sc_hd__nand2_1 _6658_ (.A(_2918_),
    .B(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__nor2_1 _6659_ (.A(_2913_),
    .B(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__nand2_1 _6660_ (.A(_2921_),
    .B(_2787_),
    .Y(_2922_));
 sky130_fd_sc_hd__nand2_1 _6661_ (.A(_2912_),
    .B(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__inv_2 _6662_ (.A(_2922_),
    .Y(_2924_));
 sky130_fd_sc_hd__nand3_1 _6663_ (.A(_2910_),
    .B(_2911_),
    .C(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__nand2_1 _6664_ (.A(_2923_),
    .B(_2925_),
    .Y(_2926_));
 sky130_fd_sc_hd__nand2_1 _6665_ (.A(_2926_),
    .B(_2747_),
    .Y(_2927_));
 sky130_fd_sc_hd__nand3_1 _6666_ (.A(_2858_),
    .B(_2904_),
    .C(_2885_),
    .Y(_2928_));
 sky130_fd_sc_hd__nand2_1 _6667_ (.A(_2928_),
    .B(_2924_),
    .Y(_2929_));
 sky130_fd_sc_hd__o21ai_1 _6668_ (.A1(_2921_),
    .A2(_2903_),
    .B1(_2787_),
    .Y(_2930_));
 sky130_fd_sc_hd__nand2_1 _6669_ (.A(_2930_),
    .B(_2889_),
    .Y(_2931_));
 sky130_fd_sc_hd__nand2_1 _6670_ (.A(_2929_),
    .B(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__nand2_1 _6671_ (.A(_2932_),
    .B(_2739_),
    .Y(_2933_));
 sky130_fd_sc_hd__nand3_1 _6672_ (.A(_2927_),
    .B(_2933_),
    .C(_2750_),
    .Y(_2934_));
 sky130_fd_sc_hd__nand2_1 _6673_ (.A(_2903_),
    .B(_2821_),
    .Y(_2935_));
 sky130_fd_sc_hd__nand2_1 _6674_ (.A(_2934_),
    .B(_2935_),
    .Y(net27));
 sky130_fd_sc_hd__or2_1 _6675_ (.A(_2916_),
    .B(_2915_),
    .X(_2936_));
 sky130_fd_sc_hd__nand2_1 _6676_ (.A(_2936_),
    .B(_2727_),
    .Y(_2937_));
 sky130_fd_sc_hd__inv_2 _6677_ (.A(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__nand2_1 _6678_ (.A(_2938_),
    .B(_2787_),
    .Y(_2939_));
 sky130_fd_sc_hd__inv_2 _6679_ (.A(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__nand2_1 _6680_ (.A(_2931_),
    .B(_2940_),
    .Y(_2941_));
 sky130_fd_sc_hd__nand3_1 _6681_ (.A(_2930_),
    .B(_2889_),
    .C(_2939_),
    .Y(_2942_));
 sky130_fd_sc_hd__nand2_1 _6682_ (.A(_2941_),
    .B(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__nand2_1 _6683_ (.A(_2943_),
    .B(_2739_),
    .Y(_2944_));
 sky130_fd_sc_hd__nand3_1 _6684_ (.A(_2925_),
    .B(_2747_),
    .C(_2939_),
    .Y(_2945_));
 sky130_fd_sc_hd__nand3_1 _6685_ (.A(_2944_),
    .B(_2750_),
    .C(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__a2111o_1 _6686_ (.A1(net18),
    .A2(_2746_),
    .B1(_3031_),
    .C1(_2913_),
    .D1(_2920_),
    .X(_2947_));
 sky130_fd_sc_hd__nand2_1 _6687_ (.A(_2946_),
    .B(_2947_),
    .Y(net28));
 sky130_fd_sc_hd__a211o_1 _6688_ (.A1(net18),
    .A2(_2746_),
    .B1(_3031_),
    .C1(_2937_),
    .X(_2948_));
 sky130_fd_sc_hd__o31ai_2 _6689_ (.A1(_2738_),
    .A2(_2741_),
    .A3(_2751_),
    .B1(_2948_),
    .Y(net29));
 sky130_fd_sc_hd__buf_4 _6690_ (.A(net19),
    .X(_2949_));
 sky130_fd_sc_hd__clkbuf_8 _6691_ (.A(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__buf_4 _6692_ (.A(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__buf_4 _6693_ (.A(net21),
    .X(_2952_));
 sky130_fd_sc_hd__clkbuf_8 _6694_ (.A(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__buf_4 _6695_ (.A(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__or2b_2 _6696_ (.A(wb_clk_i),
    .B_N(_2952_),
    .X(_2955_));
 sky130_fd_sc_hd__buf_1 _6697_ (.A(_2955_),
    .X(_2956_));
 sky130_fd_sc_hd__buf_1 _6698_ (.A(clknet_1_0__leaf__2956_),
    .X(_2957_));
 sky130_fd_sc_hd__buf_1 _6699_ (.A(clknet_1_0__leaf__2957_),
    .X(_2958_));
 sky130_fd_sc_hd__o21ai_2 _6700_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_0__leaf__2958_),
    .Y(_0000_));
 sky130_fd_sc_hd__o21ai_2 _6701_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_0__leaf__2958_),
    .Y(_0001_));
 sky130_fd_sc_hd__o21ai_2 _6702_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_0__leaf__2958_),
    .Y(_0002_));
 sky130_fd_sc_hd__o21ai_2 _6703_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_0__leaf__2958_),
    .Y(_0003_));
 sky130_fd_sc_hd__o21ai_2 _6704_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_1__leaf__2958_),
    .Y(_0004_));
 sky130_fd_sc_hd__o21ai_2 _6705_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_1__leaf__2958_),
    .Y(_0005_));
 sky130_fd_sc_hd__o21ai_2 _6706_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_1__leaf__2958_),
    .Y(_0006_));
 sky130_fd_sc_hd__o21ai_2 _6707_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_1__leaf__2958_),
    .Y(_0007_));
 sky130_fd_sc_hd__o21ai_2 _6708_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_1__leaf__2958_),
    .Y(_0008_));
 sky130_fd_sc_hd__o21ai_2 _6709_ (.A1(_2951_),
    .A2(_2954_),
    .B1(clknet_1_1__leaf__2958_),
    .Y(_0009_));
 sky130_fd_sc_hd__buf_6 _6710_ (.A(_2950_),
    .X(_2959_));
 sky130_fd_sc_hd__clkbuf_8 _6711_ (.A(_2953_),
    .X(_2960_));
 sky130_fd_sc_hd__buf_1 _6712_ (.A(clknet_1_0__leaf__2957_),
    .X(_2961_));
 sky130_fd_sc_hd__o21ai_2 _6713_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_1__leaf__2961_),
    .Y(_0010_));
 sky130_fd_sc_hd__o21ai_2 _6714_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_1__leaf__2961_),
    .Y(_0011_));
 sky130_fd_sc_hd__o21ai_2 _6715_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_1__leaf__2961_),
    .Y(_0012_));
 sky130_fd_sc_hd__o21ai_2 _6716_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_1__leaf__2961_),
    .Y(_0013_));
 sky130_fd_sc_hd__o21ai_2 _6717_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_1__leaf__2961_),
    .Y(_0014_));
 sky130_fd_sc_hd__o21ai_2 _6718_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_1__leaf__2961_),
    .Y(_0015_));
 sky130_fd_sc_hd__o21ai_2 _6719_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_0__leaf__2961_),
    .Y(_0016_));
 sky130_fd_sc_hd__o21ai_2 _6720_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_0__leaf__2961_),
    .Y(_0017_));
 sky130_fd_sc_hd__o21ai_2 _6721_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_0__leaf__2961_),
    .Y(_0018_));
 sky130_fd_sc_hd__o21ai_2 _6722_ (.A1(_2959_),
    .A2(_2960_),
    .B1(clknet_1_0__leaf__2961_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_4 _6723_ (.A(_2950_),
    .X(_2962_));
 sky130_fd_sc_hd__buf_4 _6724_ (.A(_2953_),
    .X(_2963_));
 sky130_fd_sc_hd__buf_1 _6725_ (.A(clknet_1_0__leaf__2957_),
    .X(_2964_));
 sky130_fd_sc_hd__o21ai_2 _6726_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_0__leaf__2964_),
    .Y(_0020_));
 sky130_fd_sc_hd__o21ai_2 _6727_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_0__leaf__2964_),
    .Y(_0021_));
 sky130_fd_sc_hd__o21ai_2 _6728_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_0__leaf__2964_),
    .Y(_0022_));
 sky130_fd_sc_hd__o21ai_2 _6729_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_1__leaf__2964_),
    .Y(_0023_));
 sky130_fd_sc_hd__o21ai_2 _6730_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_0__leaf__2964_),
    .Y(_0024_));
 sky130_fd_sc_hd__o21ai_2 _6731_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_1__leaf__2964_),
    .Y(_0025_));
 sky130_fd_sc_hd__o21ai_2 _6732_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_1__leaf__2964_),
    .Y(_0026_));
 sky130_fd_sc_hd__o21ai_2 _6733_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_1__leaf__2964_),
    .Y(_0027_));
 sky130_fd_sc_hd__o21ai_2 _6734_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_1__leaf__2964_),
    .Y(_0028_));
 sky130_fd_sc_hd__o21ai_2 _6735_ (.A1(_2962_),
    .A2(_2963_),
    .B1(clknet_1_1__leaf__2964_),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_4 _6736_ (.A(_2950_),
    .X(_2965_));
 sky130_fd_sc_hd__buf_4 _6737_ (.A(_2953_),
    .X(_2966_));
 sky130_fd_sc_hd__buf_1 _6738_ (.A(clknet_1_0__leaf__2957_),
    .X(_2967_));
 sky130_fd_sc_hd__o21ai_2 _6739_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_0__leaf__2967_),
    .Y(_0030_));
 sky130_fd_sc_hd__o21ai_2 _6740_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_0__leaf__2967_),
    .Y(_0031_));
 sky130_fd_sc_hd__o21ai_2 _6741_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_0__leaf__2967_),
    .Y(_0032_));
 sky130_fd_sc_hd__o21ai_2 _6742_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_0__leaf__2967_),
    .Y(_0033_));
 sky130_fd_sc_hd__o21ai_2 _6743_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_1__leaf__2967_),
    .Y(_0034_));
 sky130_fd_sc_hd__o21ai_2 _6744_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_1__leaf__2967_),
    .Y(_0035_));
 sky130_fd_sc_hd__o21ai_2 _6745_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_1__leaf__2967_),
    .Y(_0036_));
 sky130_fd_sc_hd__o21ai_2 _6746_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_1__leaf__2967_),
    .Y(_0037_));
 sky130_fd_sc_hd__o21ai_2 _6747_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_1__leaf__2967_),
    .Y(_0038_));
 sky130_fd_sc_hd__o21ai_2 _6748_ (.A1(_2965_),
    .A2(_2966_),
    .B1(clknet_1_1__leaf__2967_),
    .Y(_0039_));
 sky130_fd_sc_hd__buf_4 _6749_ (.A(_2950_),
    .X(_2968_));
 sky130_fd_sc_hd__buf_4 _6750_ (.A(_2953_),
    .X(_2969_));
 sky130_fd_sc_hd__buf_1 _6751_ (.A(clknet_1_1__leaf__2957_),
    .X(_2970_));
 sky130_fd_sc_hd__o21ai_2 _6752_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_0__leaf__2970_),
    .Y(_0040_));
 sky130_fd_sc_hd__o21ai_2 _6753_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_0__leaf__2970_),
    .Y(_0041_));
 sky130_fd_sc_hd__o21ai_2 _6754_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_0__leaf__2970_),
    .Y(_0042_));
 sky130_fd_sc_hd__o21ai_2 _6755_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_0__leaf__2970_),
    .Y(_0043_));
 sky130_fd_sc_hd__o21ai_2 _6756_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_1__leaf__2970_),
    .Y(_0044_));
 sky130_fd_sc_hd__o21ai_2 _6757_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_1__leaf__2970_),
    .Y(_0045_));
 sky130_fd_sc_hd__o21ai_2 _6758_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_1__leaf__2970_),
    .Y(_0046_));
 sky130_fd_sc_hd__o21ai_2 _6759_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_1__leaf__2970_),
    .Y(_0047_));
 sky130_fd_sc_hd__o21ai_2 _6760_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_1__leaf__2970_),
    .Y(_0048_));
 sky130_fd_sc_hd__o21ai_2 _6761_ (.A1(_2968_),
    .A2(_2969_),
    .B1(clknet_1_1__leaf__2970_),
    .Y(_0049_));
 sky130_fd_sc_hd__buf_4 _6762_ (.A(_2950_),
    .X(_2971_));
 sky130_fd_sc_hd__buf_4 _6763_ (.A(_2953_),
    .X(_2972_));
 sky130_fd_sc_hd__buf_1 _6764_ (.A(clknet_1_1__leaf__2957_),
    .X(_2973_));
 sky130_fd_sc_hd__o21ai_2 _6765_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_0__leaf__2973_),
    .Y(_0050_));
 sky130_fd_sc_hd__o21ai_2 _6766_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_0__leaf__2973_),
    .Y(_0051_));
 sky130_fd_sc_hd__o21ai_2 _6767_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_0__leaf__2973_),
    .Y(_0052_));
 sky130_fd_sc_hd__o21ai_2 _6768_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_0__leaf__2973_),
    .Y(_0053_));
 sky130_fd_sc_hd__o21ai_2 _6769_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_0__leaf__2973_),
    .Y(_0054_));
 sky130_fd_sc_hd__o21ai_2 _6770_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_0__leaf__2973_),
    .Y(_0055_));
 sky130_fd_sc_hd__o21ai_2 _6771_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_1__leaf__2973_),
    .Y(_0056_));
 sky130_fd_sc_hd__o21ai_2 _6772_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_1__leaf__2973_),
    .Y(_0057_));
 sky130_fd_sc_hd__o21ai_2 _6773_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_1__leaf__2973_),
    .Y(_0058_));
 sky130_fd_sc_hd__o21ai_2 _6774_ (.A1(_2971_),
    .A2(_2972_),
    .B1(clknet_1_1__leaf__2973_),
    .Y(_0059_));
 sky130_fd_sc_hd__buf_4 _6775_ (.A(_2950_),
    .X(_2974_));
 sky130_fd_sc_hd__buf_4 _6776_ (.A(_2953_),
    .X(_2975_));
 sky130_fd_sc_hd__buf_1 _6777_ (.A(clknet_1_1__leaf__2957_),
    .X(_2976_));
 sky130_fd_sc_hd__o21ai_2 _6778_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_1__leaf__2976_),
    .Y(_0060_));
 sky130_fd_sc_hd__o21ai_2 _6779_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_1__leaf__2976_),
    .Y(_0061_));
 sky130_fd_sc_hd__o21ai_2 _6780_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_1__leaf__2976_),
    .Y(_0062_));
 sky130_fd_sc_hd__o21ai_2 _6781_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_1__leaf__2976_),
    .Y(_0063_));
 sky130_fd_sc_hd__o21ai_2 _6782_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_1__leaf__2976_),
    .Y(_0064_));
 sky130_fd_sc_hd__o21ai_2 _6783_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_0__leaf__2976_),
    .Y(_0065_));
 sky130_fd_sc_hd__o21ai_2 _6784_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_0__leaf__2976_),
    .Y(_0066_));
 sky130_fd_sc_hd__o21ai_2 _6785_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_0__leaf__2976_),
    .Y(_0067_));
 sky130_fd_sc_hd__o21ai_2 _6786_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_0__leaf__2976_),
    .Y(_0068_));
 sky130_fd_sc_hd__o21ai_2 _6787_ (.A1(_2974_),
    .A2(_2975_),
    .B1(clknet_1_0__leaf__2976_),
    .Y(_0069_));
 sky130_fd_sc_hd__buf_4 _6788_ (.A(_2950_),
    .X(_2977_));
 sky130_fd_sc_hd__buf_4 _6789_ (.A(_2953_),
    .X(_2978_));
 sky130_fd_sc_hd__buf_1 _6790_ (.A(clknet_1_1__leaf__2957_),
    .X(_2979_));
 sky130_fd_sc_hd__o21ai_2 _6791_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_1__leaf__2979_),
    .Y(_0070_));
 sky130_fd_sc_hd__o21ai_2 _6792_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_1__leaf__2979_),
    .Y(_0071_));
 sky130_fd_sc_hd__o21ai_2 _6793_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_1__leaf__2979_),
    .Y(_0072_));
 sky130_fd_sc_hd__o21ai_2 _6794_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_1__leaf__2979_),
    .Y(_0073_));
 sky130_fd_sc_hd__o21ai_2 _6795_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_1__leaf__2979_),
    .Y(_0074_));
 sky130_fd_sc_hd__o21ai_2 _6796_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_1__leaf__2979_),
    .Y(_0075_));
 sky130_fd_sc_hd__o21ai_2 _6797_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_0__leaf__2979_),
    .Y(_0076_));
 sky130_fd_sc_hd__o21ai_2 _6798_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_0__leaf__2979_),
    .Y(_0077_));
 sky130_fd_sc_hd__o21ai_2 _6799_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_0__leaf__2979_),
    .Y(_0078_));
 sky130_fd_sc_hd__o21ai_2 _6800_ (.A1(_2977_),
    .A2(_2978_),
    .B1(clknet_1_0__leaf__2979_),
    .Y(_0079_));
 sky130_fd_sc_hd__buf_4 _6801_ (.A(_2950_),
    .X(_2980_));
 sky130_fd_sc_hd__buf_4 _6802_ (.A(_2953_),
    .X(_2981_));
 sky130_fd_sc_hd__buf_1 _6803_ (.A(clknet_1_1__leaf__2957_),
    .X(_2982_));
 sky130_fd_sc_hd__o21ai_2 _6804_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_1__leaf__2982_),
    .Y(_0080_));
 sky130_fd_sc_hd__o21ai_2 _6805_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_1__leaf__2982_),
    .Y(_0081_));
 sky130_fd_sc_hd__o21ai_2 _6806_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_1__leaf__2982_),
    .Y(_0082_));
 sky130_fd_sc_hd__o21ai_2 _6807_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_1__leaf__2982_),
    .Y(_0083_));
 sky130_fd_sc_hd__o21ai_2 _6808_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_1__leaf__2982_),
    .Y(_0084_));
 sky130_fd_sc_hd__o21ai_2 _6809_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_0__leaf__2982_),
    .Y(_0085_));
 sky130_fd_sc_hd__o21ai_2 _6810_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_0__leaf__2982_),
    .Y(_0086_));
 sky130_fd_sc_hd__o21ai_2 _6811_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_0__leaf__2982_),
    .Y(_0087_));
 sky130_fd_sc_hd__o21ai_2 _6812_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_0__leaf__2982_),
    .Y(_0088_));
 sky130_fd_sc_hd__o21ai_2 _6813_ (.A1(_2980_),
    .A2(_2981_),
    .B1(clknet_1_0__leaf__2982_),
    .Y(_0089_));
 sky130_fd_sc_hd__buf_4 _6814_ (.A(_2949_),
    .X(_2983_));
 sky130_fd_sc_hd__buf_4 _6815_ (.A(_2952_),
    .X(_2984_));
 sky130_fd_sc_hd__buf_1 _6816_ (.A(clknet_1_1__leaf__2956_),
    .X(_2985_));
 sky130_fd_sc_hd__o21ai_2 _6817_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_1__leaf__2985_),
    .Y(_0090_));
 sky130_fd_sc_hd__o21ai_2 _6818_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_1__leaf__2985_),
    .Y(_0091_));
 sky130_fd_sc_hd__o21ai_2 _6819_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_1__leaf__2985_),
    .Y(_0092_));
 sky130_fd_sc_hd__o21ai_2 _6820_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_1__leaf__2985_),
    .Y(_0093_));
 sky130_fd_sc_hd__o21ai_2 _6821_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_0__leaf__2985_),
    .Y(_0094_));
 sky130_fd_sc_hd__o21ai_2 _6822_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_0__leaf__2985_),
    .Y(_0095_));
 sky130_fd_sc_hd__o21ai_2 _6823_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_1__leaf__2985_),
    .Y(_0096_));
 sky130_fd_sc_hd__o21ai_2 _6824_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_0__leaf__2985_),
    .Y(_0097_));
 sky130_fd_sc_hd__o21ai_2 _6825_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_0__leaf__2985_),
    .Y(_0098_));
 sky130_fd_sc_hd__o21ai_2 _6826_ (.A1(_2983_),
    .A2(_2984_),
    .B1(clknet_1_0__leaf__2985_),
    .Y(_0099_));
 sky130_fd_sc_hd__buf_4 _6827_ (.A(_2949_),
    .X(_2986_));
 sky130_fd_sc_hd__buf_4 _6828_ (.A(_2952_),
    .X(_2987_));
 sky130_fd_sc_hd__buf_1 _6829_ (.A(clknet_1_1__leaf__2956_),
    .X(_2988_));
 sky130_fd_sc_hd__o21ai_2 _6830_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_0__leaf__2988_),
    .Y(_0100_));
 sky130_fd_sc_hd__o21ai_2 _6831_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_1__leaf__2988_),
    .Y(_0101_));
 sky130_fd_sc_hd__o21ai_2 _6832_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_1__leaf__2988_),
    .Y(_0102_));
 sky130_fd_sc_hd__o21ai_2 _6833_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_1__leaf__2988_),
    .Y(_0103_));
 sky130_fd_sc_hd__o21ai_2 _6834_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_1__leaf__2988_),
    .Y(_0104_));
 sky130_fd_sc_hd__o21ai_2 _6835_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_1__leaf__2988_),
    .Y(_0105_));
 sky130_fd_sc_hd__o21ai_2 _6836_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_0__leaf__2988_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ai_2 _6837_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_0__leaf__2988_),
    .Y(_0107_));
 sky130_fd_sc_hd__o21ai_2 _6838_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_1__leaf__2988_),
    .Y(_0108_));
 sky130_fd_sc_hd__o21ai_2 _6839_ (.A1(_2986_),
    .A2(_2987_),
    .B1(clknet_1_0__leaf__2988_),
    .Y(_0109_));
 sky130_fd_sc_hd__buf_4 _6840_ (.A(_2949_),
    .X(_2989_));
 sky130_fd_sc_hd__buf_4 _6841_ (.A(_2952_),
    .X(_2990_));
 sky130_fd_sc_hd__buf_1 _6842_ (.A(clknet_1_1__leaf__2956_),
    .X(_2991_));
 sky130_fd_sc_hd__o21ai_2 _6843_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_1__leaf__2991_),
    .Y(_0110_));
 sky130_fd_sc_hd__o21ai_2 _6844_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_1__leaf__2991_),
    .Y(_0111_));
 sky130_fd_sc_hd__o21ai_2 _6845_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_1__leaf__2991_),
    .Y(_0112_));
 sky130_fd_sc_hd__o21ai_2 _6846_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_1__leaf__2991_),
    .Y(_0113_));
 sky130_fd_sc_hd__o21ai_2 _6847_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_1__leaf__2991_),
    .Y(_0114_));
 sky130_fd_sc_hd__o21ai_2 _6848_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_0__leaf__2991_),
    .Y(_0115_));
 sky130_fd_sc_hd__o21ai_2 _6849_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_0__leaf__2991_),
    .Y(_0116_));
 sky130_fd_sc_hd__o21ai_2 _6850_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_0__leaf__2991_),
    .Y(_0117_));
 sky130_fd_sc_hd__o21ai_2 _6851_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_0__leaf__2991_),
    .Y(_0118_));
 sky130_fd_sc_hd__o21ai_2 _6852_ (.A1(_2989_),
    .A2(_2990_),
    .B1(clknet_1_0__leaf__2991_),
    .Y(_0119_));
 sky130_fd_sc_hd__buf_4 _6853_ (.A(_2949_),
    .X(_2992_));
 sky130_fd_sc_hd__buf_4 _6854_ (.A(_2952_),
    .X(_2993_));
 sky130_fd_sc_hd__buf_1 _6855_ (.A(clknet_1_0__leaf__2956_),
    .X(_2994_));
 sky130_fd_sc_hd__o21ai_2 _6856_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_0__leaf__2994_),
    .Y(_0120_));
 sky130_fd_sc_hd__o21ai_2 _6857_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_0__leaf__2994_),
    .Y(_0121_));
 sky130_fd_sc_hd__o21ai_2 _6858_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_0__leaf__2994_),
    .Y(_0122_));
 sky130_fd_sc_hd__o21ai_2 _6859_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_1__leaf__2994_),
    .Y(_0123_));
 sky130_fd_sc_hd__o21ai_2 _6860_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_1__leaf__2994_),
    .Y(_0124_));
 sky130_fd_sc_hd__o21ai_2 _6861_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_0__leaf__2994_),
    .Y(_0125_));
 sky130_fd_sc_hd__o21ai_2 _6862_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_1__leaf__2994_),
    .Y(_0126_));
 sky130_fd_sc_hd__o21ai_2 _6863_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_1__leaf__2994_),
    .Y(_0127_));
 sky130_fd_sc_hd__o21ai_2 _6864_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_1__leaf__2994_),
    .Y(_0128_));
 sky130_fd_sc_hd__o21ai_2 _6865_ (.A1(_2992_),
    .A2(_2993_),
    .B1(clknet_1_1__leaf__2994_),
    .Y(_0129_));
 sky130_fd_sc_hd__buf_4 _6866_ (.A(_2949_),
    .X(_2995_));
 sky130_fd_sc_hd__buf_4 _6867_ (.A(_2952_),
    .X(_2996_));
 sky130_fd_sc_hd__buf_1 _6868_ (.A(clknet_1_1__leaf__2956_),
    .X(_2997_));
 sky130_fd_sc_hd__o21ai_2 _6869_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_0__leaf__2997_),
    .Y(_0130_));
 sky130_fd_sc_hd__o21ai_2 _6870_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_1__leaf__2997_),
    .Y(_0131_));
 sky130_fd_sc_hd__o21ai_2 _6871_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_0__leaf__2997_),
    .Y(_0132_));
 sky130_fd_sc_hd__o21ai_2 _6872_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_0__leaf__2997_),
    .Y(_0133_));
 sky130_fd_sc_hd__o21ai_2 _6873_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_0__leaf__2997_),
    .Y(_0134_));
 sky130_fd_sc_hd__o21ai_2 _6874_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_0__leaf__2997_),
    .Y(_0135_));
 sky130_fd_sc_hd__o21ai_2 _6875_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_0__leaf__2997_),
    .Y(_0136_));
 sky130_fd_sc_hd__o21ai_2 _6876_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_1__leaf__2997_),
    .Y(_0137_));
 sky130_fd_sc_hd__o21ai_2 _6877_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_1__leaf__2997_),
    .Y(_0138_));
 sky130_fd_sc_hd__o21ai_2 _6878_ (.A1(_2995_),
    .A2(_2996_),
    .B1(clknet_1_1__leaf__2997_),
    .Y(_0139_));
 sky130_fd_sc_hd__buf_4 _6879_ (.A(_2949_),
    .X(_2998_));
 sky130_fd_sc_hd__buf_4 _6880_ (.A(_2952_),
    .X(_2999_));
 sky130_fd_sc_hd__buf_1 _6881_ (.A(clknet_1_0__leaf__2956_),
    .X(_3000_));
 sky130_fd_sc_hd__o21ai_2 _6882_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_1__leaf__3000_),
    .Y(_0140_));
 sky130_fd_sc_hd__o21ai_2 _6883_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_1__leaf__3000_),
    .Y(_0141_));
 sky130_fd_sc_hd__o21ai_2 _6884_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_1__leaf__3000_),
    .Y(_0142_));
 sky130_fd_sc_hd__o21ai_2 _6885_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_1__leaf__3000_),
    .Y(_0143_));
 sky130_fd_sc_hd__o21ai_2 _6886_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_1__leaf__3000_),
    .Y(_0144_));
 sky130_fd_sc_hd__o21ai_2 _6887_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_1__leaf__3000_),
    .Y(_0145_));
 sky130_fd_sc_hd__o21ai_2 _6888_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_0__leaf__3000_),
    .Y(_0146_));
 sky130_fd_sc_hd__o21ai_2 _6889_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_0__leaf__3000_),
    .Y(_0147_));
 sky130_fd_sc_hd__o21ai_2 _6890_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_0__leaf__3000_),
    .Y(_0148_));
 sky130_fd_sc_hd__o21ai_2 _6891_ (.A1(_2998_),
    .A2(_2999_),
    .B1(clknet_1_0__leaf__3000_),
    .Y(_0149_));
 sky130_fd_sc_hd__buf_4 _6892_ (.A(_2949_),
    .X(_3001_));
 sky130_fd_sc_hd__buf_4 _6893_ (.A(_2952_),
    .X(_3002_));
 sky130_fd_sc_hd__buf_1 _6894_ (.A(clknet_1_0__leaf__2956_),
    .X(_3003_));
 sky130_fd_sc_hd__o21ai_2 _6895_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_1__leaf__3003_),
    .Y(_0150_));
 sky130_fd_sc_hd__o21ai_2 _6896_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_1__leaf__3003_),
    .Y(_0151_));
 sky130_fd_sc_hd__o21ai_2 _6897_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_1__leaf__3003_),
    .Y(_0152_));
 sky130_fd_sc_hd__o21ai_2 _6898_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_1__leaf__3003_),
    .Y(_0153_));
 sky130_fd_sc_hd__o21ai_2 _6899_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_1__leaf__3003_),
    .Y(_0154_));
 sky130_fd_sc_hd__o21ai_2 _6900_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_0__leaf__3003_),
    .Y(_0155_));
 sky130_fd_sc_hd__o21ai_2 _6901_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_0__leaf__3003_),
    .Y(_0156_));
 sky130_fd_sc_hd__o21ai_2 _6902_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_0__leaf__3003_),
    .Y(_0157_));
 sky130_fd_sc_hd__o21ai_2 _6903_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_1__leaf__3003_),
    .Y(_0158_));
 sky130_fd_sc_hd__o21ai_2 _6904_ (.A1(_3001_),
    .A2(_3002_),
    .B1(clknet_1_0__leaf__3003_),
    .Y(_0159_));
 sky130_fd_sc_hd__o21ai_2 _6905_ (.A1(_2950_),
    .A2(_2953_),
    .B1(clknet_1_0__leaf__2957_),
    .Y(_0160_));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(_0000_),
    .D(_0161_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(_0001_),
    .D(_0162_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(_0002_),
    .D(_0163_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfxtp_1 _6909_ (.CLK(_0003_),
    .D(_0164_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfxtp_1 _6910_ (.CLK(_0004_),
    .D(_0165_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfxtp_1 _6911_ (.CLK(_0005_),
    .D(_0166_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfxtp_1 _6912_ (.CLK(_0006_),
    .D(_0167_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfxtp_1 _6913_ (.CLK(_0007_),
    .D(_0168_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfxtp_1 _6914_ (.CLK(_0008_),
    .D(_0169_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfxtp_1 _6915_ (.CLK(_0009_),
    .D(_0170_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfxtp_1 _6916_ (.CLK(_0010_),
    .D(_0171_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfxtp_1 _6917_ (.CLK(_0011_),
    .D(_0172_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfxtp_1 _6918_ (.CLK(_0012_),
    .D(_0173_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfxtp_1 _6919_ (.CLK(_0013_),
    .D(_0174_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfxtp_1 _6920_ (.CLK(_0014_),
    .D(_0175_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfxtp_1 _6921_ (.CLK(_0015_),
    .D(_0176_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_1 _6922_ (.CLK(_0016_),
    .D(_0177_),
    .Q(\egd_top.BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6923_ (.CLK(_0017_),
    .D(_0178_),
    .Q(\egd_top.BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6924_ (.CLK(_0018_),
    .D(_0179_),
    .Q(\egd_top.BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6925_ (.CLK(_0019_),
    .D(_0180_),
    .Q(\egd_top.BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6926_ (.CLK(_0020_),
    .D(_0181_),
    .Q(\egd_top.BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6927_ (.CLK(_0021_),
    .D(_0182_),
    .Q(\egd_top.BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6928_ (.CLK(_0022_),
    .D(_0183_),
    .Q(\egd_top.BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6929_ (.CLK(_0023_),
    .D(_0184_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfxtp_2 _6930_ (.CLK(_0024_),
    .D(_0185_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfxtp_2 _6931_ (.CLK(_0025_),
    .D(_0186_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfxtp_2 _6932_ (.CLK(_0026_),
    .D(_0187_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfxtp_1 _6933_ (.CLK(_0027_),
    .D(_0188_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfxtp_1 _6934_ (.CLK(_0028_),
    .D(_0189_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfxtp_1 _6935_ (.CLK(_0029_),
    .D(_0190_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfxtp_1 _6936_ (.CLK(_0030_),
    .D(_0191_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfxtp_1 _6937_ (.CLK(_0031_),
    .D(_0192_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfxtp_1 _6938_ (.CLK(_0032_),
    .D(_0193_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfxtp_1 _6939_ (.CLK(_0033_),
    .D(_0194_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfxtp_1 _6940_ (.CLK(_0034_),
    .D(_0195_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfxtp_1 _6941_ (.CLK(_0035_),
    .D(_0196_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfxtp_1 _6942_ (.CLK(_0036_),
    .D(_0197_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfxtp_1 _6943_ (.CLK(_0037_),
    .D(_0198_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfxtp_1 _6944_ (.CLK(_0038_),
    .D(_0199_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfxtp_1 _6945_ (.CLK(_0039_),
    .D(_0200_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfxtp_1 _6946_ (.CLK(_0040_),
    .D(_0201_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfxtp_1 _6947_ (.CLK(_0041_),
    .D(_0202_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfxtp_1 _6948_ (.CLK(_0042_),
    .D(_0203_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfxtp_1 _6949_ (.CLK(_0043_),
    .D(_0204_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfxtp_1 _6950_ (.CLK(_0044_),
    .D(_0205_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfxtp_1 _6951_ (.CLK(_0045_),
    .D(_0206_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _6952_ (.CLK(_0046_),
    .D(_0207_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _6953_ (.CLK(_0047_),
    .D(_0208_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _6954_ (.CLK(_0048_),
    .D(_0209_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _6955_ (.CLK(_0049_),
    .D(_0210_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _6956_ (.CLK(_0050_),
    .D(_0211_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _6957_ (.CLK(_0051_),
    .D(_0212_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _6958_ (.CLK(_0052_),
    .D(_0213_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _6959_ (.CLK(_0053_),
    .D(_0214_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _6960_ (.CLK(_0054_),
    .D(_0215_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _6961_ (.CLK(_0055_),
    .D(_0216_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _6962_ (.CLK(_0056_),
    .D(_0217_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _6963_ (.CLK(_0057_),
    .D(_0218_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _6964_ (.CLK(_0058_),
    .D(_0219_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _6965_ (.CLK(_0059_),
    .D(_0220_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _6966_ (.CLK(_0060_),
    .D(_0221_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _6967_ (.CLK(_0061_),
    .D(_0222_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _6968_ (.CLK(_0062_),
    .D(_0223_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _6969_ (.CLK(_0063_),
    .D(_0224_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _6970_ (.CLK(_0064_),
    .D(_0225_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _6971_ (.CLK(_0065_),
    .D(_0226_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _6972_ (.CLK(_0066_),
    .D(_0227_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _6973_ (.CLK(_0067_),
    .D(_0228_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _6974_ (.CLK(_0068_),
    .D(_0229_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(_0069_),
    .D(_0230_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(_0070_),
    .D(_0231_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(_0071_),
    .D(_0232_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(_0072_),
    .D(_0233_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(_0073_),
    .D(_0234_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _6980_ (.CLK(_0074_),
    .D(_0235_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(_0075_),
    .D(_0236_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _6982_ (.CLK(_0076_),
    .D(_0237_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(_0077_),
    .D(_0238_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(_0078_),
    .D(_0239_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(_0079_),
    .D(_0240_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _6986_ (.CLK(_0080_),
    .D(_0241_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(_0081_),
    .D(_0242_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _6988_ (.CLK(_0082_),
    .D(_0243_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(_0083_),
    .D(_0244_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _6990_ (.CLK(_0084_),
    .D(_0245_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _6991_ (.CLK(_0085_),
    .D(_0246_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _6992_ (.CLK(_0086_),
    .D(_0247_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6993_ (.CLK(_0087_),
    .D(_0248_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6994_ (.CLK(_0088_),
    .D(_0249_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6995_ (.CLK(_0089_),
    .D(_0250_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(_0090_),
    .D(_0251_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6997_ (.CLK(_0091_),
    .D(_0252_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6998_ (.CLK(_0092_),
    .D(_0253_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6999_ (.CLK(_0093_),
    .D(_0254_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7000_ (.CLK(_0094_),
    .D(_0255_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7001_ (.CLK(_0095_),
    .D(_0256_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7002_ (.CLK(_0096_),
    .D(_0257_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7003_ (.CLK(_0097_),
    .D(_0258_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7004_ (.CLK(_0098_),
    .D(_0259_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7005_ (.CLK(_0099_),
    .D(_0260_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7006_ (.CLK(_0100_),
    .D(_0261_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7007_ (.CLK(_0101_),
    .D(_0262_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_2 _7008_ (.CLK(_0102_),
    .D(_0263_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_2 _7009_ (.CLK(_0103_),
    .D(_0264_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_2 _7010_ (.CLK(_0104_),
    .D(_0265_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _7011_ (.CLK(_0105_),
    .D(_0266_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _7012_ (.CLK(_0106_),
    .D(_0267_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _7013_ (.CLK(_0107_),
    .D(_0268_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _7014_ (.CLK(_0108_),
    .D(_0269_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _7015_ (.CLK(_0109_),
    .D(_0270_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _7016_ (.CLK(_0110_),
    .D(_0271_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _7017_ (.CLK(_0111_),
    .D(_0272_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7018_ (.CLK(_0112_),
    .D(_0273_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7019_ (.CLK(_0113_),
    .D(_0274_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7020_ (.CLK(_0114_),
    .D(_0275_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7021_ (.CLK(_0115_),
    .D(_0276_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7022_ (.CLK(_0116_),
    .D(_0277_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7023_ (.CLK(_0117_),
    .D(_0278_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7024_ (.CLK(_0118_),
    .D(_0279_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7025_ (.CLK(_0119_),
    .D(_0280_),
    .Q(\egd_top.BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7026_ (.CLK(_0120_),
    .D(_0281_),
    .Q(\egd_top.BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7027_ (.CLK(_0121_),
    .D(_0282_),
    .Q(\egd_top.BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7028_ (.CLK(_0122_),
    .D(_0283_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7029_ (.CLK(_0123_),
    .D(_0284_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7030_ (.CLK(_0124_),
    .D(_0285_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7031_ (.CLK(_0125_),
    .D(_0286_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7032_ (.CLK(_0126_),
    .D(_0287_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7033_ (.CLK(_0127_),
    .D(_0288_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7034_ (.CLK(_0128_),
    .D(_0289_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7035_ (.CLK(_0129_),
    .D(_0290_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfxtp_2 _7036_ (.CLK(_0130_),
    .D(_0291_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7037_ (.CLK(_0131_),
    .D(_0292_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _7038_ (.CLK(_0132_),
    .D(_0293_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7039_ (.CLK(_0133_),
    .D(_0294_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfxtp_2 _7040_ (.CLK(_0134_),
    .D(_0295_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7041_ (.CLK(_0135_),
    .D(_0296_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7042_ (.CLK(_0136_),
    .D(_0297_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7043_ (.CLK(_0137_),
    .D(_0298_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfxtp_1 _7044_ (.CLK(_0138_),
    .D(_0299_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfxtp_1 _7045_ (.CLK(_0139_),
    .D(_0300_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfxtp_1 _7046_ (.CLK(_0140_),
    .D(_0301_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfxtp_1 _7047_ (.CLK(_0141_),
    .D(_0302_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfxtp_1 _7048_ (.CLK(_0142_),
    .D(_0303_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfxtp_1 _7049_ (.CLK(_0143_),
    .D(_0304_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfxtp_1 _7050_ (.CLK(_0144_),
    .D(_0305_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfxtp_1 _7051_ (.CLK(_0145_),
    .D(_0306_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfxtp_1 _7052_ (.CLK(_0146_),
    .D(_0307_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfxtp_1 _7053_ (.CLK(_0147_),
    .D(_0308_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfxtp_1 _7054_ (.CLK(_0148_),
    .D(_0309_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfxtp_1 _7055_ (.CLK(_0149_),
    .D(_0310_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfxtp_1 _7056_ (.CLK(_0150_),
    .D(_0311_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfxtp_1 _7057_ (.CLK(_0151_),
    .D(_0312_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfxtp_1 _7058_ (.CLK(_0152_),
    .D(_0313_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfxtp_2 _7059_ (.CLK(_0153_),
    .D(_0314_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfxtp_2 _7060_ (.CLK(_0154_),
    .D(_0315_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_2 _7061_ (.CLK(_0155_),
    .D(_0316_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_2 _7062_ (.CLK(_0156_),
    .D(_0317_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _7063_ (.CLK(_0157_),
    .D(_0318_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _7064_ (.CLK(_0158_),
    .D(_0319_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _7065_ (.CLK(_0159_),
    .D(_0320_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_2 _7066_ (.CLK(_0160_),
    .D(_0321_),
    .Q(net36));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2956_ (.A(_2956_),
    .X(clknet_0__2956_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2957_ (.A(_2957_),
    .X(clknet_0__2957_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2958_ (.A(_2958_),
    .X(clknet_0__2958_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2961_ (.A(_2961_),
    .X(clknet_0__2961_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2964_ (.A(_2964_),
    .X(clknet_0__2964_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2967_ (.A(_2967_),
    .X(clknet_0__2967_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2970_ (.A(_2970_),
    .X(clknet_0__2970_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2973_ (.A(_2973_),
    .X(clknet_0__2973_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2976_ (.A(_2976_),
    .X(clknet_0__2976_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2979_ (.A(_2979_),
    .X(clknet_0__2979_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2982_ (.A(_2982_),
    .X(clknet_0__2982_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2985_ (.A(_2985_),
    .X(clknet_0__2985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2988_ (.A(_2988_),
    .X(clknet_0__2988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2991_ (.A(_2991_),
    .X(clknet_0__2991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2994_ (.A(_2994_),
    .X(clknet_0__2994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2997_ (.A(_2997_),
    .X(clknet_0__2997_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3000_ (.A(_3000_),
    .X(clknet_0__3000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3003_ (.A(_3003_),
    .X(clknet_0__3003_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2956_ (.A(clknet_0__2956_),
    .X(clknet_1_0__leaf__2956_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2957_ (.A(clknet_0__2957_),
    .X(clknet_1_0__leaf__2957_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2958_ (.A(clknet_0__2958_),
    .X(clknet_1_0__leaf__2958_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2961_ (.A(clknet_0__2961_),
    .X(clknet_1_0__leaf__2961_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2964_ (.A(clknet_0__2964_),
    .X(clknet_1_0__leaf__2964_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2967_ (.A(clknet_0__2967_),
    .X(clknet_1_0__leaf__2967_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2970_ (.A(clknet_0__2970_),
    .X(clknet_1_0__leaf__2970_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2973_ (.A(clknet_0__2973_),
    .X(clknet_1_0__leaf__2973_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2976_ (.A(clknet_0__2976_),
    .X(clknet_1_0__leaf__2976_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2979_ (.A(clknet_0__2979_),
    .X(clknet_1_0__leaf__2979_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2982_ (.A(clknet_0__2982_),
    .X(clknet_1_0__leaf__2982_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2985_ (.A(clknet_0__2985_),
    .X(clknet_1_0__leaf__2985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2988_ (.A(clknet_0__2988_),
    .X(clknet_1_0__leaf__2988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2991_ (.A(clknet_0__2991_),
    .X(clknet_1_0__leaf__2991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2994_ (.A(clknet_0__2994_),
    .X(clknet_1_0__leaf__2994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2997_ (.A(clknet_0__2997_),
    .X(clknet_1_0__leaf__2997_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3000_ (.A(clknet_0__3000_),
    .X(clknet_1_0__leaf__3000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3003_ (.A(clknet_0__3003_),
    .X(clknet_1_0__leaf__3003_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2956_ (.A(clknet_0__2956_),
    .X(clknet_1_1__leaf__2956_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2957_ (.A(clknet_0__2957_),
    .X(clknet_1_1__leaf__2957_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2958_ (.A(clknet_0__2958_),
    .X(clknet_1_1__leaf__2958_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2961_ (.A(clknet_0__2961_),
    .X(clknet_1_1__leaf__2961_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2964_ (.A(clknet_0__2964_),
    .X(clknet_1_1__leaf__2964_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2967_ (.A(clknet_0__2967_),
    .X(clknet_1_1__leaf__2967_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2970_ (.A(clknet_0__2970_),
    .X(clknet_1_1__leaf__2970_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2973_ (.A(clknet_0__2973_),
    .X(clknet_1_1__leaf__2973_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2976_ (.A(clknet_0__2976_),
    .X(clknet_1_1__leaf__2976_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2979_ (.A(clknet_0__2979_),
    .X(clknet_1_1__leaf__2979_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2982_ (.A(clknet_0__2982_),
    .X(clknet_1_1__leaf__2982_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2985_ (.A(clknet_0__2985_),
    .X(clknet_1_1__leaf__2985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2988_ (.A(clknet_0__2988_),
    .X(clknet_1_1__leaf__2988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2991_ (.A(clknet_0__2991_),
    .X(clknet_1_1__leaf__2991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2994_ (.A(clknet_0__2994_),
    .X(clknet_1_1__leaf__2994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2997_ (.A(clknet_0__2997_),
    .X(clknet_1_1__leaf__2997_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3000_ (.A(clknet_0__3000_),
    .X(clknet_1_1__leaf__3000_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3003_ (.A(clknet_0__3003_),
    .X(clknet_1_1__leaf__3003_));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1 (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_3047_),
    .X(net38));
 sky130_fd_sc_hd__buf_1 hold3 (.A(\egd_top.BitStream_buffer.buffer_index[5] ),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_2630_),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input1 (.A(la_data_in_47_32[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(la_data_in_47_32[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(la_data_in_47_32[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(la_data_in_47_32[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(la_data_in_47_32[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(la_data_in_47_32[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(la_data_in_47_32[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(la_data_in_47_32[9]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(la_data_in_49_48[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(la_data_in_49_48[1]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(la_data_in_64),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(la_data_in_47_32[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(la_data_in_65),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(la_oenb_64),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input3 (.A(la_data_in_47_32[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(la_data_in_47_32[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(la_data_in_47_32[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(la_data_in_47_32[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(la_data_in_47_32[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(la_data_in_47_32[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(la_data_in_47_32[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(la_data_out_15_8[0]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(la_data_out_15_8[1]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(la_data_out_15_8[2]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(la_data_out_15_8[3]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(la_data_out_15_8[4]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_data_out_15_8[5]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(la_data_out_15_8[6]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(la_data_out_15_8[7]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(la_data_out_18_16[0]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(la_data_out_18_16[1]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(la_data_out_18_16[2]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(la_data_out_22_19[0]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(la_data_out_22_19[1]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(la_data_out_22_19[2]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(la_data_out_22_19[3]));
endmodule

