magic
tech sky130A
magscale 1 2
timestamp 1695953156
<< obsli1 >>
rect 1104 2159 50876 51697
<< obsm1 >>
rect 1104 1368 50876 51728
<< metal2 >>
rect 1766 0 1822 800
rect 3146 0 3202 800
rect 4526 0 4582 800
rect 5906 0 5962 800
rect 7286 0 7342 800
rect 8666 0 8722 800
rect 10046 0 10102 800
rect 11426 0 11482 800
rect 12806 0 12862 800
rect 14186 0 14242 800
rect 15566 0 15622 800
rect 16946 0 17002 800
rect 18326 0 18382 800
rect 19706 0 19762 800
rect 21086 0 21142 800
rect 22466 0 22522 800
rect 23846 0 23902 800
rect 25226 0 25282 800
rect 26606 0 26662 800
rect 27986 0 28042 800
rect 29366 0 29422 800
rect 30746 0 30802 800
rect 32126 0 32182 800
rect 33506 0 33562 800
rect 34886 0 34942 800
rect 36266 0 36322 800
rect 37646 0 37702 800
rect 39026 0 39082 800
rect 40406 0 40462 800
rect 41786 0 41842 800
rect 43166 0 43222 800
rect 44546 0 44602 800
rect 45926 0 45982 800
rect 47306 0 47362 800
rect 48686 0 48742 800
rect 50066 0 50122 800
<< obsm2 >>
rect 1768 856 50856 51717
rect 1878 734 3090 856
rect 3258 734 4470 856
rect 4638 734 5850 856
rect 6018 734 7230 856
rect 7398 734 8610 856
rect 8778 734 9990 856
rect 10158 734 11370 856
rect 11538 734 12750 856
rect 12918 734 14130 856
rect 14298 734 15510 856
rect 15678 734 16890 856
rect 17058 734 18270 856
rect 18438 734 19650 856
rect 19818 734 21030 856
rect 21198 734 22410 856
rect 22578 734 23790 856
rect 23958 734 25170 856
rect 25338 734 26550 856
rect 26718 734 27930 856
rect 28098 734 29310 856
rect 29478 734 30690 856
rect 30858 734 32070 856
rect 32238 734 33450 856
rect 33618 734 34830 856
rect 34998 734 36210 856
rect 36378 734 37590 856
rect 37758 734 38970 856
rect 39138 734 40350 856
rect 40518 734 41730 856
rect 41898 734 43110 856
rect 43278 734 44490 856
rect 44658 734 45870 856
rect 46038 734 47250 856
rect 47418 734 48630 856
rect 48798 734 50010 856
rect 50178 734 50856 856
<< metal3 >>
rect 0 26936 800 27056
<< obsm3 >>
rect 800 27136 50771 51713
rect 880 26856 50771 27136
rect 800 1939 50771 26856
<< metal4 >>
rect 4208 2128 4528 51728
rect 19568 2128 19888 51728
rect 34928 2128 35248 51728
rect 50288 2128 50608 51728
<< obsm4 >>
rect 9259 2075 19488 44301
rect 19968 2075 34848 44301
rect 35328 2075 48885 44301
<< labels >>
rlabel metal2 s 22466 0 22522 800 6 la_data_in_47_32[0]
port 1 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in_47_32[10]
port 2 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_data_in_47_32[11]
port 3 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in_47_32[12]
port 4 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in_47_32[13]
port 5 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_data_in_47_32[14]
port 6 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in_47_32[15]
port 7 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_data_in_47_32[1]
port 8 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_data_in_47_32[2]
port 9 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_data_in_47_32[3]
port 10 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_data_in_47_32[4]
port 11 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_data_in_47_32[5]
port 12 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_data_in_47_32[6]
port 13 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_data_in_47_32[7]
port 14 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_data_in_47_32[8]
port 15 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_data_in_47_32[9]
port 16 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_data_in_49_48[0]
port 17 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in_49_48[1]
port 18 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in_64
port 19 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in_65
port 20 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 la_data_out_15_8[0]
port 21 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 la_data_out_15_8[1]
port 22 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 la_data_out_15_8[2]
port 23 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 la_data_out_15_8[3]
port 24 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 la_data_out_15_8[4]
port 25 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 la_data_out_15_8[5]
port 26 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 la_data_out_15_8[6]
port 27 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 la_data_out_15_8[7]
port 28 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 la_data_out_18_16[0]
port 29 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 la_data_out_18_16[1]
port 30 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 la_data_out_18_16[2]
port 31 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 la_data_out_22_19[0]
port 32 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 la_data_out_22_19[1]
port 33 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 la_data_out_22_19[2]
port 34 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 la_data_out_22_19[3]
port 35 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_oenb_64
port 36 nsew signal input
rlabel metal4 s 4208 2128 4528 51728 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 51728 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 51728 6 vssd1
port 38 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 51728 6 vssd1
port 38 nsew ground bidirectional
rlabel metal3 s 0 26936 800 27056 6 wb_clk_i
port 39 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 51995 54139
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9903962
string GDS_FILE /home/uniccass/H.264_Decoder/openlane/egd_top_wrapper/runs/23_09_28_18_32/results/signoff/egd_top_wrapper.magic.gds
string GDS_START 551578
<< end >>

