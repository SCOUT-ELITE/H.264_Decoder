// This is the unpowered netlist.
module egd_top_wrapper (la_data_in_64,
    la_data_in_65,
    la_oenb_64,
    la_oenb_65,
    wb_clk_i,
    wb_rst_i,
    la_data_in_47_32,
    la_data_in_49_48,
    la_data_out_15_8,
    la_data_out_18_16,
    la_data_out_22_19);
 input la_data_in_64;
 input la_data_in_65;
 input la_oenb_64;
 input la_oenb_65;
 input wb_clk_i;
 input wb_rst_i;
 input [15:0] la_data_in_47_32;
 input [1:0] la_data_in_49_48;
 output [7:0] la_data_out_15_8;
 output [2:0] la_data_out_18_16;
 output [3:0] la_data_out_22_19;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire clknet_0__3030_;
 wire clknet_0__3031_;
 wire clknet_0__3032_;
 wire clknet_0__3035_;
 wire clknet_0__3038_;
 wire clknet_0__3041_;
 wire clknet_0__3044_;
 wire clknet_0__3047_;
 wire clknet_0__3050_;
 wire clknet_0__3053_;
 wire clknet_0__3056_;
 wire clknet_0__3059_;
 wire clknet_0__3062_;
 wire clknet_0__3065_;
 wire clknet_0__3068_;
 wire clknet_0__3071_;
 wire clknet_0__3074_;
 wire clknet_0__3077_;
 wire clknet_1_0__leaf__3030_;
 wire clknet_1_0__leaf__3031_;
 wire clknet_1_0__leaf__3032_;
 wire clknet_1_0__leaf__3035_;
 wire clknet_1_0__leaf__3038_;
 wire clknet_1_0__leaf__3041_;
 wire clknet_1_0__leaf__3044_;
 wire clknet_1_0__leaf__3047_;
 wire clknet_1_0__leaf__3050_;
 wire clknet_1_0__leaf__3053_;
 wire clknet_1_0__leaf__3056_;
 wire clknet_1_0__leaf__3059_;
 wire clknet_1_0__leaf__3062_;
 wire clknet_1_0__leaf__3065_;
 wire clknet_1_0__leaf__3068_;
 wire clknet_1_0__leaf__3071_;
 wire clknet_1_0__leaf__3074_;
 wire clknet_1_0__leaf__3077_;
 wire clknet_1_1__leaf__3030_;
 wire clknet_1_1__leaf__3031_;
 wire clknet_1_1__leaf__3032_;
 wire clknet_1_1__leaf__3035_;
 wire clknet_1_1__leaf__3038_;
 wire clknet_1_1__leaf__3041_;
 wire clknet_1_1__leaf__3044_;
 wire clknet_1_1__leaf__3047_;
 wire clknet_1_1__leaf__3050_;
 wire clknet_1_1__leaf__3053_;
 wire clknet_1_1__leaf__3056_;
 wire clknet_1_1__leaf__3059_;
 wire clknet_1_1__leaf__3062_;
 wire clknet_1_1__leaf__3065_;
 wire clknet_1_1__leaf__3068_;
 wire clknet_1_1__leaf__3071_;
 wire clknet_1_1__leaf__3074_;
 wire clknet_1_1__leaf__3077_;
 wire \egd_top.BitStream_buffer.BS_buffer[0] ;
 wire \egd_top.BitStream_buffer.BS_buffer[100] ;
 wire \egd_top.BitStream_buffer.BS_buffer[101] ;
 wire \egd_top.BitStream_buffer.BS_buffer[102] ;
 wire \egd_top.BitStream_buffer.BS_buffer[103] ;
 wire \egd_top.BitStream_buffer.BS_buffer[104] ;
 wire \egd_top.BitStream_buffer.BS_buffer[105] ;
 wire \egd_top.BitStream_buffer.BS_buffer[106] ;
 wire \egd_top.BitStream_buffer.BS_buffer[107] ;
 wire \egd_top.BitStream_buffer.BS_buffer[108] ;
 wire \egd_top.BitStream_buffer.BS_buffer[109] ;
 wire \egd_top.BitStream_buffer.BS_buffer[10] ;
 wire \egd_top.BitStream_buffer.BS_buffer[110] ;
 wire \egd_top.BitStream_buffer.BS_buffer[111] ;
 wire \egd_top.BitStream_buffer.BS_buffer[112] ;
 wire \egd_top.BitStream_buffer.BS_buffer[113] ;
 wire \egd_top.BitStream_buffer.BS_buffer[114] ;
 wire \egd_top.BitStream_buffer.BS_buffer[115] ;
 wire \egd_top.BitStream_buffer.BS_buffer[116] ;
 wire \egd_top.BitStream_buffer.BS_buffer[117] ;
 wire \egd_top.BitStream_buffer.BS_buffer[118] ;
 wire \egd_top.BitStream_buffer.BS_buffer[119] ;
 wire \egd_top.BitStream_buffer.BS_buffer[11] ;
 wire \egd_top.BitStream_buffer.BS_buffer[120] ;
 wire \egd_top.BitStream_buffer.BS_buffer[121] ;
 wire \egd_top.BitStream_buffer.BS_buffer[122] ;
 wire \egd_top.BitStream_buffer.BS_buffer[123] ;
 wire \egd_top.BitStream_buffer.BS_buffer[124] ;
 wire \egd_top.BitStream_buffer.BS_buffer[125] ;
 wire \egd_top.BitStream_buffer.BS_buffer[126] ;
 wire \egd_top.BitStream_buffer.BS_buffer[127] ;
 wire \egd_top.BitStream_buffer.BS_buffer[12] ;
 wire \egd_top.BitStream_buffer.BS_buffer[13] ;
 wire \egd_top.BitStream_buffer.BS_buffer[14] ;
 wire \egd_top.BitStream_buffer.BS_buffer[15] ;
 wire \egd_top.BitStream_buffer.BS_buffer[16] ;
 wire \egd_top.BitStream_buffer.BS_buffer[17] ;
 wire \egd_top.BitStream_buffer.BS_buffer[18] ;
 wire \egd_top.BitStream_buffer.BS_buffer[19] ;
 wire \egd_top.BitStream_buffer.BS_buffer[1] ;
 wire \egd_top.BitStream_buffer.BS_buffer[20] ;
 wire \egd_top.BitStream_buffer.BS_buffer[21] ;
 wire \egd_top.BitStream_buffer.BS_buffer[22] ;
 wire \egd_top.BitStream_buffer.BS_buffer[23] ;
 wire \egd_top.BitStream_buffer.BS_buffer[24] ;
 wire \egd_top.BitStream_buffer.BS_buffer[25] ;
 wire \egd_top.BitStream_buffer.BS_buffer[26] ;
 wire \egd_top.BitStream_buffer.BS_buffer[27] ;
 wire \egd_top.BitStream_buffer.BS_buffer[28] ;
 wire \egd_top.BitStream_buffer.BS_buffer[29] ;
 wire \egd_top.BitStream_buffer.BS_buffer[2] ;
 wire \egd_top.BitStream_buffer.BS_buffer[30] ;
 wire \egd_top.BitStream_buffer.BS_buffer[31] ;
 wire \egd_top.BitStream_buffer.BS_buffer[32] ;
 wire \egd_top.BitStream_buffer.BS_buffer[33] ;
 wire \egd_top.BitStream_buffer.BS_buffer[34] ;
 wire \egd_top.BitStream_buffer.BS_buffer[35] ;
 wire \egd_top.BitStream_buffer.BS_buffer[36] ;
 wire \egd_top.BitStream_buffer.BS_buffer[37] ;
 wire \egd_top.BitStream_buffer.BS_buffer[38] ;
 wire \egd_top.BitStream_buffer.BS_buffer[39] ;
 wire \egd_top.BitStream_buffer.BS_buffer[3] ;
 wire \egd_top.BitStream_buffer.BS_buffer[40] ;
 wire \egd_top.BitStream_buffer.BS_buffer[41] ;
 wire \egd_top.BitStream_buffer.BS_buffer[42] ;
 wire \egd_top.BitStream_buffer.BS_buffer[43] ;
 wire \egd_top.BitStream_buffer.BS_buffer[44] ;
 wire \egd_top.BitStream_buffer.BS_buffer[45] ;
 wire \egd_top.BitStream_buffer.BS_buffer[46] ;
 wire \egd_top.BitStream_buffer.BS_buffer[47] ;
 wire \egd_top.BitStream_buffer.BS_buffer[48] ;
 wire \egd_top.BitStream_buffer.BS_buffer[49] ;
 wire \egd_top.BitStream_buffer.BS_buffer[4] ;
 wire \egd_top.BitStream_buffer.BS_buffer[50] ;
 wire \egd_top.BitStream_buffer.BS_buffer[51] ;
 wire \egd_top.BitStream_buffer.BS_buffer[52] ;
 wire \egd_top.BitStream_buffer.BS_buffer[53] ;
 wire \egd_top.BitStream_buffer.BS_buffer[54] ;
 wire \egd_top.BitStream_buffer.BS_buffer[55] ;
 wire \egd_top.BitStream_buffer.BS_buffer[56] ;
 wire \egd_top.BitStream_buffer.BS_buffer[57] ;
 wire \egd_top.BitStream_buffer.BS_buffer[58] ;
 wire \egd_top.BitStream_buffer.BS_buffer[59] ;
 wire \egd_top.BitStream_buffer.BS_buffer[5] ;
 wire \egd_top.BitStream_buffer.BS_buffer[60] ;
 wire \egd_top.BitStream_buffer.BS_buffer[61] ;
 wire \egd_top.BitStream_buffer.BS_buffer[62] ;
 wire \egd_top.BitStream_buffer.BS_buffer[63] ;
 wire \egd_top.BitStream_buffer.BS_buffer[64] ;
 wire \egd_top.BitStream_buffer.BS_buffer[65] ;
 wire \egd_top.BitStream_buffer.BS_buffer[66] ;
 wire \egd_top.BitStream_buffer.BS_buffer[67] ;
 wire \egd_top.BitStream_buffer.BS_buffer[68] ;
 wire \egd_top.BitStream_buffer.BS_buffer[69] ;
 wire \egd_top.BitStream_buffer.BS_buffer[6] ;
 wire \egd_top.BitStream_buffer.BS_buffer[70] ;
 wire \egd_top.BitStream_buffer.BS_buffer[71] ;
 wire \egd_top.BitStream_buffer.BS_buffer[72] ;
 wire \egd_top.BitStream_buffer.BS_buffer[73] ;
 wire \egd_top.BitStream_buffer.BS_buffer[74] ;
 wire \egd_top.BitStream_buffer.BS_buffer[75] ;
 wire \egd_top.BitStream_buffer.BS_buffer[76] ;
 wire \egd_top.BitStream_buffer.BS_buffer[77] ;
 wire \egd_top.BitStream_buffer.BS_buffer[78] ;
 wire \egd_top.BitStream_buffer.BS_buffer[79] ;
 wire \egd_top.BitStream_buffer.BS_buffer[7] ;
 wire \egd_top.BitStream_buffer.BS_buffer[80] ;
 wire \egd_top.BitStream_buffer.BS_buffer[81] ;
 wire \egd_top.BitStream_buffer.BS_buffer[82] ;
 wire \egd_top.BitStream_buffer.BS_buffer[83] ;
 wire \egd_top.BitStream_buffer.BS_buffer[84] ;
 wire \egd_top.BitStream_buffer.BS_buffer[85] ;
 wire \egd_top.BitStream_buffer.BS_buffer[86] ;
 wire \egd_top.BitStream_buffer.BS_buffer[87] ;
 wire \egd_top.BitStream_buffer.BS_buffer[88] ;
 wire \egd_top.BitStream_buffer.BS_buffer[89] ;
 wire \egd_top.BitStream_buffer.BS_buffer[8] ;
 wire \egd_top.BitStream_buffer.BS_buffer[90] ;
 wire \egd_top.BitStream_buffer.BS_buffer[91] ;
 wire \egd_top.BitStream_buffer.BS_buffer[92] ;
 wire \egd_top.BitStream_buffer.BS_buffer[93] ;
 wire \egd_top.BitStream_buffer.BS_buffer[94] ;
 wire \egd_top.BitStream_buffer.BS_buffer[95] ;
 wire \egd_top.BitStream_buffer.BS_buffer[96] ;
 wire \egd_top.BitStream_buffer.BS_buffer[97] ;
 wire \egd_top.BitStream_buffer.BS_buffer[98] ;
 wire \egd_top.BitStream_buffer.BS_buffer[99] ;
 wire \egd_top.BitStream_buffer.BS_buffer[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[10] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[11] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[12] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[13] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[14] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[15] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[1] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[2] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[3] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[4] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[5] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[6] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[7] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[8] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_valid_n ;
 wire \egd_top.BitStream_buffer.buffer_index[4] ;
 wire \egd_top.BitStream_buffer.buffer_index[5] ;
 wire \egd_top.BitStream_buffer.buffer_index[6] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[1] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[2] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[3] ;
 wire \egd_top.BitStream_buffer.pc[1] ;
 wire \egd_top.BitStream_buffer.pc[2] ;
 wire \egd_top.BitStream_buffer.pc[3] ;
 wire \egd_top.BitStream_buffer.pc[4] ;
 wire \egd_top.BitStream_buffer.pc[5] ;
 wire \egd_top.BitStream_buffer.pc[6] ;
 wire \egd_top.BitStream_buffer.pc_previous[0] ;
 wire \egd_top.BitStream_buffer.pc_previous[1] ;
 wire \egd_top.BitStream_buffer.pc_previous[2] ;
 wire \egd_top.BitStream_buffer.pc_previous[3] ;
 wire \egd_top.BitStream_buffer.pc_previous[4] ;
 wire \egd_top.BitStream_buffer.pc_previous[5] ;
 wire \egd_top.BitStream_buffer.pc_previous[6] ;
 wire \egd_top.exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_2282_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_3242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_3242_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_1717_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net6));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__or2b_4 _3516_ (.A(net23),
    .B_N(net22),
    .X(_3078_));
 sky130_fd_sc_hd__o21a_4 _3517_ (.A1(net20),
    .A2(net22),
    .B1(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__buf_6 _3518_ (.A(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__buf_2 _3519_ (.A(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__inv_2 _3520_ (.A(net37),
    .Y(_3082_));
 sky130_fd_sc_hd__nand2_1 _3521_ (.A(net36),
    .B(net35),
    .Y(_3083_));
 sky130_fd_sc_hd__inv_2 _3522_ (.A(net38),
    .Y(_3084_));
 sky130_fd_sc_hd__o21ai_1 _3523_ (.A1(_3082_),
    .A2(_3083_),
    .B1(_3084_),
    .Y(_3085_));
 sky130_fd_sc_hd__nand2_1 _3524_ (.A(_3081_),
    .B(_3085_),
    .Y(_3086_));
 sky130_fd_sc_hd__inv_2 _3525_ (.A(_3086_),
    .Y(_0321_));
 sky130_fd_sc_hd__a21o_1 _3526_ (.A1(_3082_),
    .A2(_3083_),
    .B1(_3085_),
    .X(_3087_));
 sky130_fd_sc_hd__nand2_1 _3527_ (.A(net38),
    .B(net37),
    .Y(_3088_));
 sky130_fd_sc_hd__inv_2 _3528_ (.A(_3079_),
    .Y(_3089_));
 sky130_fd_sc_hd__clkbuf_4 _3529_ (.A(_3089_),
    .X(_3090_));
 sky130_fd_sc_hd__a21oi_1 _3530_ (.A1(_3087_),
    .A2(_3088_),
    .B1(_3090_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _3531_ (.A(net35),
    .Y(_3091_));
 sky130_fd_sc_hd__nor2_1 _3532_ (.A(net37),
    .B(net36),
    .Y(_3092_));
 sky130_fd_sc_hd__nor2_1 _3533_ (.A(_3084_),
    .B(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__nor2_1 _3534_ (.A(_3091_),
    .B(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__or2_1 _3535_ (.A(net36),
    .B(_3094_),
    .X(_3095_));
 sky130_fd_sc_hd__nand2_1 _3536_ (.A(_3094_),
    .B(net36),
    .Y(_3096_));
 sky130_fd_sc_hd__and3_1 _3537_ (.A(_3095_),
    .B(_3080_),
    .C(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__clkbuf_1 _3538_ (.A(_3097_),
    .X(_0319_));
 sky130_fd_sc_hd__inv_2 _3539_ (.A(_3093_),
    .Y(_3098_));
 sky130_fd_sc_hd__nor2_1 _3540_ (.A(net35),
    .B(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__or3_1 _3541_ (.A(_3094_),
    .B(_3099_),
    .C(_3089_),
    .X(_3100_));
 sky130_fd_sc_hd__inv_2 _3542_ (.A(_3100_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _3543_ (.A(net34),
    .Y(_3101_));
 sky130_fd_sc_hd__nor2_1 _3544_ (.A(net33),
    .B(net32),
    .Y(_3102_));
 sky130_fd_sc_hd__nor2_1 _3545_ (.A(_3101_),
    .B(_3102_),
    .Y(_3103_));
 sky130_fd_sc_hd__a21o_1 _3546_ (.A1(net33),
    .A2(net32),
    .B1(net34),
    .X(_3104_));
 sky130_fd_sc_hd__and2b_1 _3547_ (.A_N(_3103_),
    .B(_3104_),
    .X(_3105_));
 sky130_fd_sc_hd__inv_2 _3548_ (.A(_3102_),
    .Y(_3106_));
 sky130_fd_sc_hd__nor2_1 _3549_ (.A(net34),
    .B(_3106_),
    .Y(_3107_));
 sky130_fd_sc_hd__inv_2 _3550_ (.A(_3107_),
    .Y(_3108_));
 sky130_fd_sc_hd__inv_2 _3551_ (.A(net18),
    .Y(_3109_));
 sky130_fd_sc_hd__inv_2 _3552_ (.A(net17),
    .Y(_3110_));
 sky130_fd_sc_hd__nand2_2 _3553_ (.A(_3109_),
    .B(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__or2_1 _3554_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__nand2_4 _3555_ (.A(_3111_),
    .B(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_3113_));
 sky130_fd_sc_hd__nand2_2 _3556_ (.A(_3112_),
    .B(_3113_),
    .Y(_3114_));
 sky130_fd_sc_hd__inv_2 _3557_ (.A(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__nand2_2 _3558_ (.A(_3115_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3116_));
 sky130_fd_sc_hd__inv_2 _3559_ (.A(_3116_),
    .Y(_3117_));
 sky130_fd_sc_hd__and3_1 _3560_ (.A(_3117_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3118_));
 sky130_fd_sc_hd__buf_6 _3561_ (.A(_3118_),
    .X(_3119_));
 sky130_fd_sc_hd__inv_2 _3562_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_3120_));
 sky130_fd_sc_hd__and3_2 _3563_ (.A(_3120_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3121_));
 sky130_fd_sc_hd__nand2_2 _3564_ (.A(_3119_),
    .B(_3121_),
    .Y(_3122_));
 sky130_fd_sc_hd__inv_2 _3565_ (.A(_3122_),
    .Y(_3123_));
 sky130_fd_sc_hd__inv_2 _3566_ (.A(net44),
    .Y(_3124_));
 sky130_fd_sc_hd__inv_2 _3567_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_3125_));
 sky130_fd_sc_hd__and3_1 _3568_ (.A(_3124_),
    .B(_3125_),
    .C(net47),
    .X(_3126_));
 sky130_fd_sc_hd__or4b_1 _3569_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_3108_),
    .C(_3123_),
    .D_N(_3126_),
    .X(_3127_));
 sky130_fd_sc_hd__or3b_1 _3570_ (.A(_3101_),
    .B(net33),
    .C_N(net32),
    .X(_3128_));
 sky130_fd_sc_hd__nor2_1 _3571_ (.A(_3103_),
    .B(_3107_),
    .Y(_3129_));
 sky130_fd_sc_hd__inv_2 _3572_ (.A(_3129_),
    .Y(_3130_));
 sky130_fd_sc_hd__nand3_1 _3573_ (.A(_3127_),
    .B(_3128_),
    .C(_3130_),
    .Y(_3131_));
 sky130_fd_sc_hd__inv_2 _3574_ (.A(net42),
    .Y(_3132_));
 sky130_fd_sc_hd__and3_1 _3575_ (.A(_3132_),
    .B(_3124_),
    .C(_3125_),
    .X(_3133_));
 sky130_fd_sc_hd__and4_1 _3576_ (.A(\egd_top.BitStream_buffer.pc_previous[0] ),
    .B(\egd_top.BitStream_buffer.pc_previous[1] ),
    .C(\egd_top.BitStream_buffer.pc_previous[2] ),
    .D(\egd_top.BitStream_buffer.pc_previous[3] ),
    .X(_3134_));
 sky130_fd_sc_hd__a31o_1 _3577_ (.A1(_3134_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .A3(\egd_top.BitStream_buffer.pc_previous[5] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[6] ),
    .X(_3135_));
 sky130_fd_sc_hd__or3b_1 _3578_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_3123_),
    .C_N(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__or2_1 _3579_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_3120_),
    .X(_3137_));
 sky130_fd_sc_hd__a21oi_1 _3580_ (.A1(_3136_),
    .A2(_3137_),
    .B1(_3108_),
    .Y(_3138_));
 sky130_fd_sc_hd__a31o_1 _3581_ (.A1(\egd_top.BitStream_buffer.pc[6] ),
    .A2(_3107_),
    .A3(_3133_),
    .B1(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__or2_1 _3582_ (.A(_3131_),
    .B(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__and4_1 _3583_ (.A(_3082_),
    .B(_3091_),
    .C(net38),
    .D(net36),
    .X(_3141_));
 sky130_fd_sc_hd__nand2_1 _3584_ (.A(_3140_),
    .B(_3141_),
    .Y(_3142_));
 sky130_fd_sc_hd__nand2_1 _3585_ (.A(_3142_),
    .B(_3101_),
    .Y(_3143_));
 sky130_fd_sc_hd__o211a_1 _3586_ (.A1(_3105_),
    .A2(_3142_),
    .B1(_3081_),
    .C1(_3143_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _3587_ (.A(_3102_),
    .B(_3104_),
    .Y(_3144_));
 sky130_fd_sc_hd__a21o_1 _3588_ (.A1(_3140_),
    .A2(_3141_),
    .B1(net33),
    .X(_3145_));
 sky130_fd_sc_hd__o211a_1 _3589_ (.A1(_3142_),
    .A2(_3144_),
    .B1(_3081_),
    .C1(_3145_),
    .X(_0316_));
 sky130_fd_sc_hd__o21ai_1 _3590_ (.A1(net32),
    .A2(_3130_),
    .B1(_3127_),
    .Y(_3146_));
 sky130_fd_sc_hd__o21bai_1 _3591_ (.A1(_3139_),
    .A2(_3146_),
    .B1_N(_3142_),
    .Y(_3147_));
 sky130_fd_sc_hd__nand2_1 _3592_ (.A(_3142_),
    .B(net32),
    .Y(_3148_));
 sky130_fd_sc_hd__a21oi_1 _3593_ (.A1(_3147_),
    .A2(_3148_),
    .B1(_3090_),
    .Y(_0315_));
 sky130_fd_sc_hd__buf_6 _3594_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .X(_3149_));
 sky130_fd_sc_hd__inv_2 _3595_ (.A(_3149_),
    .Y(_3150_));
 sky130_fd_sc_hd__clkbuf_4 _3596_ (.A(_3150_),
    .X(_3151_));
 sky130_fd_sc_hd__o21ai_1 _3597_ (.A1(_3151_),
    .A2(_3141_),
    .B1(_3081_),
    .Y(_0314_));
 sky130_fd_sc_hd__buf_2 _3598_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .X(_3152_));
 sky130_fd_sc_hd__or2_1 _3599_ (.A(net34),
    .B(net33),
    .X(_3153_));
 sky130_fd_sc_hd__nand2_1 _3600_ (.A(net34),
    .B(net33),
    .Y(_3154_));
 sky130_fd_sc_hd__nand2_1 _3601_ (.A(_3092_),
    .B(_3084_),
    .Y(_3155_));
 sky130_fd_sc_hd__a22o_2 _3602_ (.A1(_3153_),
    .A2(_3154_),
    .B1(_3098_),
    .B2(_3155_),
    .X(_3156_));
 sky130_fd_sc_hd__or4b_2 _3603_ (.A(_3132_),
    .B(_3124_),
    .C(_3125_),
    .D_N(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__buf_2 _3604_ (.A(_3157_),
    .X(_3158_));
 sky130_fd_sc_hd__clkbuf_4 _3605_ (.A(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__mux2_1 _3606_ (.A0(net7),
    .A1(_3152_),
    .S(_3159_),
    .X(_3160_));
 sky130_fd_sc_hd__buf_6 _3607_ (.A(_3080_),
    .X(_3161_));
 sky130_fd_sc_hd__and2_1 _3608_ (.A(_3160_),
    .B(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__clkbuf_1 _3609_ (.A(_3162_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_4 _3610_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_3163_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(net6),
    .A1(_3163_),
    .S(_3159_),
    .X(_3164_));
 sky130_fd_sc_hd__buf_8 _3612_ (.A(_3079_),
    .X(_3165_));
 sky130_fd_sc_hd__buf_6 _3613_ (.A(_3165_),
    .X(_3166_));
 sky130_fd_sc_hd__and2_1 _3614_ (.A(_3164_),
    .B(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__clkbuf_1 _3615_ (.A(_3167_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_2 _3616_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .X(_3168_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(net5),
    .A1(_3168_),
    .S(_3159_),
    .X(_3169_));
 sky130_fd_sc_hd__and2_1 _3618_ (.A(_3169_),
    .B(_3166_),
    .X(_3170_));
 sky130_fd_sc_hd__clkbuf_1 _3619_ (.A(_3170_),
    .X(_0311_));
 sky130_fd_sc_hd__buf_2 _3620_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .X(_3171_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(net4),
    .A1(_3171_),
    .S(_3159_),
    .X(_3172_));
 sky130_fd_sc_hd__and2_1 _3622_ (.A(_3172_),
    .B(_3166_),
    .X(_3173_));
 sky130_fd_sc_hd__clkbuf_1 _3623_ (.A(_3173_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_4 _3624_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .X(_3174_));
 sky130_fd_sc_hd__mux2_1 _3625_ (.A0(net3),
    .A1(_3174_),
    .S(_3159_),
    .X(_3175_));
 sky130_fd_sc_hd__and2_1 _3626_ (.A(_3175_),
    .B(_3166_),
    .X(_3176_));
 sky130_fd_sc_hd__clkbuf_1 _3627_ (.A(_3176_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_2 _3628_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .X(_3177_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(net2),
    .A1(_3177_),
    .S(_3159_),
    .X(_3178_));
 sky130_fd_sc_hd__and2_1 _3630_ (.A(_3178_),
    .B(_3166_),
    .X(_3179_));
 sky130_fd_sc_hd__clkbuf_1 _3631_ (.A(_3179_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_2 _3632_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .X(_3180_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(net16),
    .A1(_3180_),
    .S(_3159_),
    .X(_3181_));
 sky130_fd_sc_hd__and2_4 _3634_ (.A(_3181_),
    .B(_3166_),
    .X(_3182_));
 sky130_fd_sc_hd__clkbuf_1 _3635_ (.A(_3182_),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_4 _3636_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_3183_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(net15),
    .A1(_3183_),
    .S(_3159_),
    .X(_3184_));
 sky130_fd_sc_hd__and2_1 _3638_ (.A(_3184_),
    .B(_3166_),
    .X(_3185_));
 sky130_fd_sc_hd__clkbuf_1 _3639_ (.A(_3185_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_2 _3640_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_3186_));
 sky130_fd_sc_hd__mux2_1 _3641_ (.A0(net14),
    .A1(_3186_),
    .S(_3159_),
    .X(_3187_));
 sky130_fd_sc_hd__and2_1 _3642_ (.A(_3187_),
    .B(_3166_),
    .X(_3188_));
 sky130_fd_sc_hd__clkbuf_1 _3643_ (.A(_3188_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_2 _3644_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_3189_));
 sky130_fd_sc_hd__mux2_1 _3645_ (.A0(net13),
    .A1(_3189_),
    .S(_3159_),
    .X(_3190_));
 sky130_fd_sc_hd__and2_1 _3646_ (.A(_3190_),
    .B(_3166_),
    .X(_3191_));
 sky130_fd_sc_hd__clkbuf_1 _3647_ (.A(_3191_),
    .X(_0304_));
 sky130_fd_sc_hd__buf_2 _3648_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_3192_));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(net12),
    .A1(_3192_),
    .S(_3158_),
    .X(_3193_));
 sky130_fd_sc_hd__and2_4 _3650_ (.A(_3193_),
    .B(_3166_),
    .X(_3194_));
 sky130_fd_sc_hd__clkbuf_1 _3651_ (.A(_3194_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_4 _3652_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .X(_3195_));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(net11),
    .A1(_3195_),
    .S(_3158_),
    .X(_3196_));
 sky130_fd_sc_hd__buf_8 _3654_ (.A(_3165_),
    .X(_3197_));
 sky130_fd_sc_hd__and2_1 _3655_ (.A(_3196_),
    .B(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__clkbuf_1 _3656_ (.A(_3198_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_2 _3657_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_3199_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(net10),
    .A1(_3199_),
    .S(_3158_),
    .X(_3200_));
 sky130_fd_sc_hd__and2_1 _3659_ (.A(_3200_),
    .B(_3197_),
    .X(_3201_));
 sky130_fd_sc_hd__clkbuf_1 _3660_ (.A(_3201_),
    .X(_0301_));
 sky130_fd_sc_hd__buf_2 _3661_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_3202_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(net9),
    .A1(_3202_),
    .S(_3158_),
    .X(_3203_));
 sky130_fd_sc_hd__and2_1 _3663_ (.A(_3203_),
    .B(_3197_),
    .X(_3204_));
 sky130_fd_sc_hd__clkbuf_1 _3664_ (.A(_3204_),
    .X(_0300_));
 sky130_fd_sc_hd__buf_2 _3665_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_3205_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(net8),
    .A1(_3205_),
    .S(_3158_),
    .X(_3206_));
 sky130_fd_sc_hd__and2_1 _3667_ (.A(_3206_),
    .B(_3197_),
    .X(_3207_));
 sky130_fd_sc_hd__clkbuf_1 _3668_ (.A(_3207_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_2 _3669_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_3208_));
 sky130_fd_sc_hd__mux2_1 _3670_ (.A0(net1),
    .A1(_3208_),
    .S(_3158_),
    .X(_3209_));
 sky130_fd_sc_hd__and2_1 _3671_ (.A(_3209_),
    .B(_3197_),
    .X(_3210_));
 sky130_fd_sc_hd__clkbuf_1 _3672_ (.A(_3210_),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_1 _3673_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B1(_3081_),
    .Y(_3211_));
 sky130_fd_sc_hd__buf_2 _3674_ (.A(_3149_),
    .X(_3212_));
 sky130_fd_sc_hd__clkbuf_4 _3675_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .X(_3213_));
 sky130_fd_sc_hd__nand2_2 _3676_ (.A(_3114_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3214_));
 sky130_fd_sc_hd__inv_2 _3677_ (.A(_3214_),
    .Y(_3215_));
 sky130_fd_sc_hd__inv_2 _3678_ (.A(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3216_));
 sky130_fd_sc_hd__and3_4 _3679_ (.A(_3215_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3216_),
    .X(_3217_));
 sky130_fd_sc_hd__inv_2 _3680_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_3218_));
 sky130_fd_sc_hd__and3_2 _3681_ (.A(_3120_),
    .B(_3218_),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_3219_));
 sky130_fd_sc_hd__buf_2 _3682_ (.A(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__and2_1 _3683_ (.A(_3217_),
    .B(_3220_),
    .X(_3221_));
 sky130_fd_sc_hd__clkbuf_2 _3684_ (.A(_3221_),
    .X(_3222_));
 sky130_fd_sc_hd__buf_2 _3685_ (.A(_3222_),
    .X(_3223_));
 sky130_fd_sc_hd__clkbuf_4 _3686_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .X(_3224_));
 sky130_fd_sc_hd__and3_1 _3687_ (.A(_3117_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3216_),
    .X(_3225_));
 sky130_fd_sc_hd__buf_4 _3688_ (.A(_3225_),
    .X(_3226_));
 sky130_fd_sc_hd__and2_1 _3689_ (.A(_3226_),
    .B(_3220_),
    .X(_3227_));
 sky130_fd_sc_hd__clkbuf_2 _3690_ (.A(_3227_),
    .X(_3228_));
 sky130_fd_sc_hd__buf_2 _3691_ (.A(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__inv_2 _3692_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_3230_));
 sky130_fd_sc_hd__nand2_2 _3693_ (.A(_3115_),
    .B(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__inv_2 _3694_ (.A(_3231_),
    .Y(_3232_));
 sky130_fd_sc_hd__and3_1 _3695_ (.A(_3232_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3216_),
    .X(_3233_));
 sky130_fd_sc_hd__clkbuf_8 _3696_ (.A(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__and2_1 _3697_ (.A(_3234_),
    .B(_3219_),
    .X(_3235_));
 sky130_fd_sc_hd__clkbuf_2 _3698_ (.A(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__buf_2 _3699_ (.A(_3236_),
    .X(_3237_));
 sky130_fd_sc_hd__clkbuf_4 _3700_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .X(_3238_));
 sky130_fd_sc_hd__nand2_1 _3701_ (.A(_3237_),
    .B(_3238_),
    .Y(_3239_));
 sky130_fd_sc_hd__nand2_4 _3702_ (.A(_3114_),
    .B(_3230_),
    .Y(_3240_));
 sky130_fd_sc_hd__inv_2 _3703_ (.A(_3240_),
    .Y(_3241_));
 sky130_fd_sc_hd__and3_4 _3704_ (.A(_3241_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_3216_),
    .X(_3242_));
 sky130_fd_sc_hd__and2_1 _3705_ (.A(_3242_),
    .B(_3219_),
    .X(_3243_));
 sky130_fd_sc_hd__clkbuf_2 _3706_ (.A(_3243_),
    .X(_3244_));
 sky130_fd_sc_hd__buf_2 _3707_ (.A(_3244_),
    .X(_3245_));
 sky130_fd_sc_hd__clkbuf_4 _3708_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .X(_3246_));
 sky130_fd_sc_hd__nand2_1 _3709_ (.A(_3245_),
    .B(_3246_),
    .Y(_3247_));
 sky130_fd_sc_hd__nand2_1 _3710_ (.A(_3239_),
    .B(_3247_),
    .Y(_3248_));
 sky130_fd_sc_hd__a221oi_1 _3711_ (.A1(_3213_),
    .A2(_3223_),
    .B1(_3224_),
    .B2(_3229_),
    .C1(_3248_),
    .Y(_3249_));
 sky130_fd_sc_hd__clkbuf_4 _3712_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_3250_));
 sky130_fd_sc_hd__and3_4 _3713_ (.A(_3215_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3251_));
 sky130_fd_sc_hd__and2_1 _3714_ (.A(_3251_),
    .B(_3220_),
    .X(_3252_));
 sky130_fd_sc_hd__clkbuf_2 _3715_ (.A(_3252_),
    .X(_3253_));
 sky130_fd_sc_hd__buf_2 _3716_ (.A(_3253_),
    .X(_3254_));
 sky130_fd_sc_hd__clkbuf_4 _3717_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_3255_));
 sky130_fd_sc_hd__and2_1 _3718_ (.A(_3119_),
    .B(_3220_),
    .X(_3256_));
 sky130_fd_sc_hd__clkbuf_2 _3719_ (.A(_3256_),
    .X(_3257_));
 sky130_fd_sc_hd__buf_2 _3720_ (.A(_3257_),
    .X(_3258_));
 sky130_fd_sc_hd__and3_1 _3721_ (.A(_3232_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3259_));
 sky130_fd_sc_hd__buf_4 _3722_ (.A(_3259_),
    .X(_3260_));
 sky130_fd_sc_hd__and2_1 _3723_ (.A(_3260_),
    .B(_3219_),
    .X(_3261_));
 sky130_fd_sc_hd__clkbuf_2 _3724_ (.A(_3261_),
    .X(_3262_));
 sky130_fd_sc_hd__buf_2 _3725_ (.A(_3262_),
    .X(_3263_));
 sky130_fd_sc_hd__clkbuf_4 _3726_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_3264_));
 sky130_fd_sc_hd__nand2_1 _3727_ (.A(_3263_),
    .B(_3264_),
    .Y(_3265_));
 sky130_fd_sc_hd__and3_1 _3728_ (.A(_3241_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_3266_));
 sky130_fd_sc_hd__buf_4 _3729_ (.A(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__and2_1 _3730_ (.A(_3267_),
    .B(_3219_),
    .X(_3268_));
 sky130_fd_sc_hd__clkbuf_2 _3731_ (.A(_3268_),
    .X(_3269_));
 sky130_fd_sc_hd__buf_2 _3732_ (.A(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_4 _3733_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_3271_));
 sky130_fd_sc_hd__nand2_1 _3734_ (.A(_3270_),
    .B(_3271_),
    .Y(_3272_));
 sky130_fd_sc_hd__nand2_1 _3735_ (.A(_3265_),
    .B(_3272_),
    .Y(_3273_));
 sky130_fd_sc_hd__a221oi_2 _3736_ (.A1(_3250_),
    .A2(_3254_),
    .B1(_3255_),
    .B2(_3258_),
    .C1(_3273_),
    .Y(_3274_));
 sky130_fd_sc_hd__clkbuf_4 _3737_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .X(_3275_));
 sky130_fd_sc_hd__inv_2 _3738_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_3276_));
 sky130_fd_sc_hd__nand2_4 _3739_ (.A(_3276_),
    .B(_3216_),
    .Y(_3277_));
 sky130_fd_sc_hd__nor2_8 _3740_ (.A(_3277_),
    .B(_3240_),
    .Y(_3278_));
 sky130_fd_sc_hd__and2_1 _3741_ (.A(_3278_),
    .B(_3220_),
    .X(_3279_));
 sky130_fd_sc_hd__clkbuf_2 _3742_ (.A(_3279_),
    .X(_3280_));
 sky130_fd_sc_hd__clkbuf_4 _3743_ (.A(_3280_),
    .X(_3281_));
 sky130_fd_sc_hd__or2_2 _3744_ (.A(_3277_),
    .B(_3231_),
    .X(_3282_));
 sky130_fd_sc_hd__inv_2 _3745_ (.A(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__and2_1 _3746_ (.A(_3283_),
    .B(_3220_),
    .X(_3284_));
 sky130_fd_sc_hd__clkbuf_2 _3747_ (.A(_3284_),
    .X(_3285_));
 sky130_fd_sc_hd__buf_2 _3748_ (.A(_3285_),
    .X(_3286_));
 sky130_fd_sc_hd__clkbuf_4 _3749_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .X(_3287_));
 sky130_fd_sc_hd__inv_2 _3750_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .Y(_3288_));
 sky130_fd_sc_hd__nor2_4 _3751_ (.A(_3277_),
    .B(_3214_),
    .Y(_3289_));
 sky130_fd_sc_hd__nand2_2 _3752_ (.A(_3289_),
    .B(_3220_),
    .Y(_3290_));
 sky130_fd_sc_hd__buf_2 _3753_ (.A(_3290_),
    .X(_3291_));
 sky130_fd_sc_hd__nor2_4 _3754_ (.A(_3277_),
    .B(_3116_),
    .Y(_3292_));
 sky130_fd_sc_hd__and2_1 _3755_ (.A(_3292_),
    .B(_3219_),
    .X(_3293_));
 sky130_fd_sc_hd__clkbuf_2 _3756_ (.A(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__buf_2 _3757_ (.A(_3294_),
    .X(_3295_));
 sky130_fd_sc_hd__clkbuf_4 _3758_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .X(_3296_));
 sky130_fd_sc_hd__nand2_1 _3759_ (.A(_3295_),
    .B(_3296_),
    .Y(_3297_));
 sky130_fd_sc_hd__o21ai_1 _3760_ (.A1(_3288_),
    .A2(_3291_),
    .B1(_3297_),
    .Y(_3298_));
 sky130_fd_sc_hd__a221oi_1 _3761_ (.A1(_3275_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_3287_),
    .C1(_3298_),
    .Y(_3299_));
 sky130_fd_sc_hd__clkbuf_4 _3762_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .X(_3300_));
 sky130_fd_sc_hd__nand2_8 _3763_ (.A(_3276_),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_3301_));
 sky130_fd_sc_hd__nor2_4 _3764_ (.A(_3301_),
    .B(_3214_),
    .Y(_3302_));
 sky130_fd_sc_hd__and2_1 _3765_ (.A(_3302_),
    .B(_3219_),
    .X(_3303_));
 sky130_fd_sc_hd__clkbuf_2 _3766_ (.A(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__buf_2 _3767_ (.A(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__clkbuf_4 _3768_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .X(_3306_));
 sky130_fd_sc_hd__nor2_4 _3769_ (.A(_3301_),
    .B(_3116_),
    .Y(_3307_));
 sky130_fd_sc_hd__and2_1 _3770_ (.A(_3307_),
    .B(_3220_),
    .X(_3308_));
 sky130_fd_sc_hd__clkbuf_2 _3771_ (.A(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__buf_2 _3772_ (.A(_3309_),
    .X(_3310_));
 sky130_fd_sc_hd__inv_2 _3773_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .Y(_3311_));
 sky130_fd_sc_hd__nor2_8 _3774_ (.A(_3301_),
    .B(_3240_),
    .Y(_3312_));
 sky130_fd_sc_hd__nand2_2 _3775_ (.A(_3312_),
    .B(_3220_),
    .Y(_3313_));
 sky130_fd_sc_hd__buf_2 _3776_ (.A(_3313_),
    .X(_3314_));
 sky130_fd_sc_hd__inv_2 _3777_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .Y(_3315_));
 sky130_fd_sc_hd__nor2_8 _3778_ (.A(_3301_),
    .B(_3231_),
    .Y(_3316_));
 sky130_fd_sc_hd__nand2_2 _3779_ (.A(_3316_),
    .B(_3220_),
    .Y(_3317_));
 sky130_fd_sc_hd__buf_2 _3780_ (.A(_3317_),
    .X(_3318_));
 sky130_fd_sc_hd__o22ai_1 _3781_ (.A1(_3311_),
    .A2(_3314_),
    .B1(_3315_),
    .B2(_3318_),
    .Y(_3319_));
 sky130_fd_sc_hd__a221oi_1 _3782_ (.A1(_3300_),
    .A2(_3305_),
    .B1(_3306_),
    .B2(_3310_),
    .C1(_3319_),
    .Y(_3320_));
 sky130_fd_sc_hd__and4_1 _3783_ (.A(_3249_),
    .B(_3274_),
    .C(_3299_),
    .D(_3320_),
    .X(_3321_));
 sky130_fd_sc_hd__clkbuf_4 _3784_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .X(_3322_));
 sky130_fd_sc_hd__buf_2 _3785_ (.A(_3121_),
    .X(_3323_));
 sky130_fd_sc_hd__and2_1 _3786_ (.A(_3267_),
    .B(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__clkbuf_2 _3787_ (.A(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__buf_2 _3788_ (.A(_3325_),
    .X(_3326_));
 sky130_fd_sc_hd__clkbuf_4 _3789_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .X(_3327_));
 sky130_fd_sc_hd__and2_1 _3790_ (.A(_3260_),
    .B(_3323_),
    .X(_3328_));
 sky130_fd_sc_hd__clkbuf_2 _3791_ (.A(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__buf_2 _3792_ (.A(_3329_),
    .X(_3330_));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_3331_));
 sky130_fd_sc_hd__clkbuf_4 _3794_ (.A(_3122_),
    .X(_3332_));
 sky130_fd_sc_hd__and2_1 _3795_ (.A(_3251_),
    .B(_3121_),
    .X(_3333_));
 sky130_fd_sc_hd__clkbuf_2 _3796_ (.A(_3333_),
    .X(_3334_));
 sky130_fd_sc_hd__buf_2 _3797_ (.A(_3334_),
    .X(_3335_));
 sky130_fd_sc_hd__clkbuf_4 _3798_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .X(_3336_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(_3335_),
    .B(_3336_),
    .Y(_3337_));
 sky130_fd_sc_hd__o21ai_1 _3800_ (.A1(_3331_),
    .A2(_3332_),
    .B1(_3337_),
    .Y(_3338_));
 sky130_fd_sc_hd__a221oi_1 _3801_ (.A1(_3322_),
    .A2(_3326_),
    .B1(_3327_),
    .B2(_3330_),
    .C1(_3338_),
    .Y(_3339_));
 sky130_fd_sc_hd__buf_2 _3802_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_3340_));
 sky130_fd_sc_hd__and2_1 _3803_ (.A(_3242_),
    .B(_3323_),
    .X(_3341_));
 sky130_fd_sc_hd__clkbuf_2 _3804_ (.A(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__buf_2 _3805_ (.A(_3342_),
    .X(_3343_));
 sky130_fd_sc_hd__clkbuf_4 _3806_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .X(_3344_));
 sky130_fd_sc_hd__and2_1 _3807_ (.A(_3234_),
    .B(_3323_),
    .X(_3345_));
 sky130_fd_sc_hd__clkbuf_2 _3808_ (.A(_3345_),
    .X(_3346_));
 sky130_fd_sc_hd__buf_2 _3809_ (.A(_3346_),
    .X(_3347_));
 sky130_fd_sc_hd__inv_2 _3810_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_3348_));
 sky130_fd_sc_hd__nand2_2 _3811_ (.A(_3226_),
    .B(_3323_),
    .Y(_3349_));
 sky130_fd_sc_hd__clkbuf_4 _3812_ (.A(_3349_),
    .X(_3350_));
 sky130_fd_sc_hd__and2_1 _3813_ (.A(_3217_),
    .B(_3121_),
    .X(_3351_));
 sky130_fd_sc_hd__clkbuf_2 _3814_ (.A(_3351_),
    .X(_3352_));
 sky130_fd_sc_hd__buf_2 _3815_ (.A(_3352_),
    .X(_3353_));
 sky130_fd_sc_hd__clkbuf_4 _3816_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .X(_3354_));
 sky130_fd_sc_hd__nand2_1 _3817_ (.A(_3353_),
    .B(_3354_),
    .Y(_3355_));
 sky130_fd_sc_hd__o21ai_1 _3818_ (.A1(_3348_),
    .A2(_3350_),
    .B1(_3355_),
    .Y(_3356_));
 sky130_fd_sc_hd__a221oi_1 _3819_ (.A1(_3340_),
    .A2(_3343_),
    .B1(_3344_),
    .B2(_3347_),
    .C1(_3356_),
    .Y(_3357_));
 sky130_fd_sc_hd__buf_2 _3820_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_3358_));
 sky130_fd_sc_hd__and2_1 _3821_ (.A(_3289_),
    .B(_3323_),
    .X(_3359_));
 sky130_fd_sc_hd__clkbuf_2 _3822_ (.A(_3359_),
    .X(_3360_));
 sky130_fd_sc_hd__buf_2 _3823_ (.A(_3360_),
    .X(_3361_));
 sky130_fd_sc_hd__buf_2 _3824_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_3362_));
 sky130_fd_sc_hd__and2_1 _3825_ (.A(_3292_),
    .B(_3323_),
    .X(_3363_));
 sky130_fd_sc_hd__clkbuf_2 _3826_ (.A(_3363_),
    .X(_3364_));
 sky130_fd_sc_hd__buf_2 _3827_ (.A(_3364_),
    .X(_3365_));
 sky130_fd_sc_hd__inv_2 _3828_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .Y(_3366_));
 sky130_fd_sc_hd__nand2_2 _3829_ (.A(_3278_),
    .B(_3323_),
    .Y(_3367_));
 sky130_fd_sc_hd__buf_2 _3830_ (.A(_3367_),
    .X(_3368_));
 sky130_fd_sc_hd__and2_1 _3831_ (.A(_3283_),
    .B(_3121_),
    .X(_3369_));
 sky130_fd_sc_hd__clkbuf_2 _3832_ (.A(_3369_),
    .X(_3370_));
 sky130_fd_sc_hd__buf_4 _3833_ (.A(_3370_),
    .X(_3371_));
 sky130_fd_sc_hd__buf_2 _3834_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_3372_));
 sky130_fd_sc_hd__nand2_1 _3835_ (.A(_3371_),
    .B(_3372_),
    .Y(_3373_));
 sky130_fd_sc_hd__o21ai_1 _3836_ (.A1(_3366_),
    .A2(_3368_),
    .B1(_3373_),
    .Y(_3374_));
 sky130_fd_sc_hd__a221oi_1 _3837_ (.A1(_3358_),
    .A2(_3361_),
    .B1(_3362_),
    .B2(_3365_),
    .C1(_3374_),
    .Y(_3375_));
 sky130_fd_sc_hd__buf_2 _3838_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .X(_3376_));
 sky130_fd_sc_hd__and2_1 _3839_ (.A(_3302_),
    .B(_3323_),
    .X(_3377_));
 sky130_fd_sc_hd__buf_2 _3840_ (.A(_3377_),
    .X(_3378_));
 sky130_fd_sc_hd__clkbuf_4 _3841_ (.A(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__buf_2 _3842_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .X(_3380_));
 sky130_fd_sc_hd__and2_1 _3843_ (.A(_3307_),
    .B(_3323_),
    .X(_3381_));
 sky130_fd_sc_hd__buf_2 _3844_ (.A(_3381_),
    .X(_3382_));
 sky130_fd_sc_hd__clkbuf_4 _3845_ (.A(_3382_),
    .X(_3383_));
 sky130_fd_sc_hd__and2_1 _3846_ (.A(_3316_),
    .B(_3121_),
    .X(_3384_));
 sky130_fd_sc_hd__clkbuf_2 _3847_ (.A(_3384_),
    .X(_3385_));
 sky130_fd_sc_hd__buf_2 _3848_ (.A(_3385_),
    .X(_3386_));
 sky130_fd_sc_hd__nand2_1 _3849_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_3387_));
 sky130_fd_sc_hd__and2_1 _3850_ (.A(_3312_),
    .B(_3121_),
    .X(_3388_));
 sky130_fd_sc_hd__clkbuf_2 _3851_ (.A(_3388_),
    .X(_3389_));
 sky130_fd_sc_hd__buf_2 _3852_ (.A(_3389_),
    .X(_3390_));
 sky130_fd_sc_hd__nand2_1 _3853_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_3391_));
 sky130_fd_sc_hd__nand2_1 _3854_ (.A(_3387_),
    .B(_3391_),
    .Y(_3392_));
 sky130_fd_sc_hd__a221oi_1 _3855_ (.A1(_3376_),
    .A2(_3379_),
    .B1(_3380_),
    .B2(_3383_),
    .C1(_3392_),
    .Y(_3393_));
 sky130_fd_sc_hd__and4_1 _3856_ (.A(_3339_),
    .B(_3357_),
    .C(_3375_),
    .D(_3393_),
    .X(_3394_));
 sky130_fd_sc_hd__clkbuf_4 _3857_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_3395_));
 sky130_fd_sc_hd__inv_2 _3858_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_3396_));
 sky130_fd_sc_hd__and3_2 _3859_ (.A(_3120_),
    .B(_3396_),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_3397_));
 sky130_fd_sc_hd__clkbuf_4 _3860_ (.A(_3397_),
    .X(_3398_));
 sky130_fd_sc_hd__and2_1 _3861_ (.A(_3217_),
    .B(_3398_),
    .X(_3399_));
 sky130_fd_sc_hd__clkbuf_2 _3862_ (.A(_3399_),
    .X(_3400_));
 sky130_fd_sc_hd__buf_2 _3863_ (.A(_3400_),
    .X(_3401_));
 sky130_fd_sc_hd__clkbuf_4 _3864_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_3402_));
 sky130_fd_sc_hd__and2_1 _3865_ (.A(_3226_),
    .B(_3398_),
    .X(_3403_));
 sky130_fd_sc_hd__clkbuf_2 _3866_ (.A(_3403_),
    .X(_3404_));
 sky130_fd_sc_hd__buf_2 _3867_ (.A(_3404_),
    .X(_3405_));
 sky130_fd_sc_hd__inv_2 _3868_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_3406_));
 sky130_fd_sc_hd__nand2_2 _3869_ (.A(_3242_),
    .B(_3398_),
    .Y(_3407_));
 sky130_fd_sc_hd__buf_2 _3870_ (.A(_3407_),
    .X(_3408_));
 sky130_fd_sc_hd__inv_2 _3871_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .Y(_3409_));
 sky130_fd_sc_hd__nand2_2 _3872_ (.A(_3234_),
    .B(_3398_),
    .Y(_3410_));
 sky130_fd_sc_hd__buf_2 _3873_ (.A(_3410_),
    .X(_3411_));
 sky130_fd_sc_hd__o22ai_1 _3874_ (.A1(_3406_),
    .A2(_3408_),
    .B1(_3409_),
    .B2(_3411_),
    .Y(_3412_));
 sky130_fd_sc_hd__a221oi_1 _3875_ (.A1(_3395_),
    .A2(_3401_),
    .B1(_3402_),
    .B2(_3405_),
    .C1(_3412_),
    .Y(_3413_));
 sky130_fd_sc_hd__buf_2 _3876_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_3414_));
 sky130_fd_sc_hd__and2_1 _3877_ (.A(_3267_),
    .B(_3398_),
    .X(_3415_));
 sky130_fd_sc_hd__clkbuf_2 _3878_ (.A(_3415_),
    .X(_3416_));
 sky130_fd_sc_hd__buf_2 _3879_ (.A(_3416_),
    .X(_3417_));
 sky130_fd_sc_hd__buf_2 _3880_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_3418_));
 sky130_fd_sc_hd__and2_1 _3881_ (.A(_3260_),
    .B(_3398_),
    .X(_3419_));
 sky130_fd_sc_hd__clkbuf_2 _3882_ (.A(_3419_),
    .X(_3420_));
 sky130_fd_sc_hd__buf_2 _3883_ (.A(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__inv_2 _3884_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_3422_));
 sky130_fd_sc_hd__nand2_2 _3885_ (.A(_3119_),
    .B(_3398_),
    .Y(_3423_));
 sky130_fd_sc_hd__buf_2 _3886_ (.A(_3423_),
    .X(_3424_));
 sky130_fd_sc_hd__and2_1 _3887_ (.A(_3251_),
    .B(_3397_),
    .X(_3425_));
 sky130_fd_sc_hd__clkbuf_2 _3888_ (.A(_3425_),
    .X(_3426_));
 sky130_fd_sc_hd__buf_2 _3889_ (.A(_3426_),
    .X(_3427_));
 sky130_fd_sc_hd__buf_2 _3890_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_3428_));
 sky130_fd_sc_hd__nand2_1 _3891_ (.A(_3427_),
    .B(_3428_),
    .Y(_3429_));
 sky130_fd_sc_hd__o21ai_1 _3892_ (.A1(_3422_),
    .A2(_3424_),
    .B1(_3429_),
    .Y(_3430_));
 sky130_fd_sc_hd__a221oi_1 _3893_ (.A1(_3414_),
    .A2(_3417_),
    .B1(_3418_),
    .B2(_3421_),
    .C1(_3430_),
    .Y(_3431_));
 sky130_fd_sc_hd__clkbuf_4 _3894_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_3432_));
 sky130_fd_sc_hd__and2_1 _3895_ (.A(_3278_),
    .B(_3397_),
    .X(_3433_));
 sky130_fd_sc_hd__clkbuf_2 _3896_ (.A(_3433_),
    .X(_3434_));
 sky130_fd_sc_hd__buf_2 _3897_ (.A(_3434_),
    .X(_3435_));
 sky130_fd_sc_hd__and2_1 _3898_ (.A(_3283_),
    .B(_3398_),
    .X(_3436_));
 sky130_fd_sc_hd__clkbuf_2 _3899_ (.A(_3436_),
    .X(_3437_));
 sky130_fd_sc_hd__buf_2 _3900_ (.A(_3437_),
    .X(_3438_));
 sky130_fd_sc_hd__clkbuf_4 _3901_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_3439_));
 sky130_fd_sc_hd__inv_2 _3902_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_3440_));
 sky130_fd_sc_hd__nand2_2 _3903_ (.A(_3289_),
    .B(_3398_),
    .Y(_3441_));
 sky130_fd_sc_hd__clkbuf_4 _3904_ (.A(_3441_),
    .X(_3442_));
 sky130_fd_sc_hd__and2_1 _3905_ (.A(_3292_),
    .B(_3397_),
    .X(_3443_));
 sky130_fd_sc_hd__clkbuf_2 _3906_ (.A(_3443_),
    .X(_3444_));
 sky130_fd_sc_hd__buf_2 _3907_ (.A(_3444_),
    .X(_3445_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_3446_));
 sky130_fd_sc_hd__o21ai_1 _3909_ (.A1(_3440_),
    .A2(_3442_),
    .B1(_3446_),
    .Y(_3447_));
 sky130_fd_sc_hd__a221oi_1 _3910_ (.A1(_3432_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_3439_),
    .C1(_3447_),
    .Y(_3448_));
 sky130_fd_sc_hd__buf_2 _3911_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_3449_));
 sky130_fd_sc_hd__and2_1 _3912_ (.A(_3302_),
    .B(_3397_),
    .X(_3450_));
 sky130_fd_sc_hd__clkbuf_2 _3913_ (.A(_3450_),
    .X(_3451_));
 sky130_fd_sc_hd__buf_2 _3914_ (.A(_3451_),
    .X(_3452_));
 sky130_fd_sc_hd__buf_2 _3915_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_3453_));
 sky130_fd_sc_hd__and2_1 _3916_ (.A(_3307_),
    .B(_3398_),
    .X(_3454_));
 sky130_fd_sc_hd__clkbuf_2 _3917_ (.A(_3454_),
    .X(_3455_));
 sky130_fd_sc_hd__buf_2 _3918_ (.A(_3455_),
    .X(_3456_));
 sky130_fd_sc_hd__and2_1 _3919_ (.A(_3316_),
    .B(_3397_),
    .X(_3457_));
 sky130_fd_sc_hd__clkbuf_2 _3920_ (.A(_3457_),
    .X(_3458_));
 sky130_fd_sc_hd__buf_2 _3921_ (.A(_3458_),
    .X(_3459_));
 sky130_fd_sc_hd__nand2_1 _3922_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_3460_));
 sky130_fd_sc_hd__and2_1 _3923_ (.A(_3312_),
    .B(_3397_),
    .X(_3461_));
 sky130_fd_sc_hd__clkbuf_2 _3924_ (.A(_3461_),
    .X(_3462_));
 sky130_fd_sc_hd__buf_4 _3925_ (.A(_3462_),
    .X(_3463_));
 sky130_fd_sc_hd__nand2_1 _3926_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_3464_));
 sky130_fd_sc_hd__nand2_1 _3927_ (.A(_3460_),
    .B(_3464_),
    .Y(_3465_));
 sky130_fd_sc_hd__a221oi_1 _3928_ (.A1(_3449_),
    .A2(_3452_),
    .B1(_3453_),
    .B2(_3456_),
    .C1(_3465_),
    .Y(_3466_));
 sky130_fd_sc_hd__and4_1 _3929_ (.A(_3413_),
    .B(_3431_),
    .C(_3448_),
    .D(_3466_),
    .X(_3467_));
 sky130_fd_sc_hd__inv_2 _3930_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .Y(_3468_));
 sky130_fd_sc_hd__and3_2 _3931_ (.A(_3120_),
    .B(_3396_),
    .C(_3218_),
    .X(_3469_));
 sky130_fd_sc_hd__buf_4 _3932_ (.A(_3469_),
    .X(_3470_));
 sky130_fd_sc_hd__nand2_2 _3933_ (.A(_3234_),
    .B(_3470_),
    .Y(_3471_));
 sky130_fd_sc_hd__buf_2 _3934_ (.A(_3471_),
    .X(_3472_));
 sky130_fd_sc_hd__and2_1 _3935_ (.A(_3217_),
    .B(_3469_),
    .X(_3473_));
 sky130_fd_sc_hd__clkbuf_2 _3936_ (.A(_3473_),
    .X(_3474_));
 sky130_fd_sc_hd__buf_2 _3937_ (.A(_3474_),
    .X(_3475_));
 sky130_fd_sc_hd__clkbuf_4 _3938_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_3476_));
 sky130_fd_sc_hd__nand2_1 _3939_ (.A(_3475_),
    .B(_3476_),
    .Y(_3477_));
 sky130_fd_sc_hd__and2_1 _3940_ (.A(_3242_),
    .B(_3469_),
    .X(_3478_));
 sky130_fd_sc_hd__clkbuf_2 _3941_ (.A(_3478_),
    .X(_3479_));
 sky130_fd_sc_hd__buf_2 _3942_ (.A(_3479_),
    .X(_3480_));
 sky130_fd_sc_hd__nand2_1 _3943_ (.A(_3480_),
    .B(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_3481_));
 sky130_fd_sc_hd__clkbuf_4 _3944_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .X(_3482_));
 sky130_fd_sc_hd__inv_2 _3945_ (.A(_3482_),
    .Y(_3483_));
 sky130_fd_sc_hd__nand2_1 _3946_ (.A(_3226_),
    .B(_3470_),
    .Y(_3484_));
 sky130_fd_sc_hd__clkbuf_2 _3947_ (.A(_3484_),
    .X(_3485_));
 sky130_fd_sc_hd__or2_1 _3948_ (.A(_3483_),
    .B(_3485_),
    .X(_3486_));
 sky130_fd_sc_hd__o2111a_1 _3949_ (.A1(_3468_),
    .A2(_3472_),
    .B1(_3477_),
    .C1(_3481_),
    .D1(_3486_),
    .X(_3487_));
 sky130_fd_sc_hd__inv_2 _3950_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .Y(_3488_));
 sky130_fd_sc_hd__nand2_2 _3951_ (.A(_3289_),
    .B(_3470_),
    .Y(_3489_));
 sky130_fd_sc_hd__buf_2 _3952_ (.A(_3489_),
    .X(_3490_));
 sky130_fd_sc_hd__inv_2 _3953_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_3491_));
 sky130_fd_sc_hd__nand2_2 _3954_ (.A(_3283_),
    .B(_3470_),
    .Y(_3492_));
 sky130_fd_sc_hd__buf_2 _3955_ (.A(_3492_),
    .X(_3493_));
 sky130_fd_sc_hd__and2_1 _3956_ (.A(_3292_),
    .B(_3470_),
    .X(_3494_));
 sky130_fd_sc_hd__clkbuf_2 _3957_ (.A(_3494_),
    .X(_3495_));
 sky130_fd_sc_hd__buf_2 _3958_ (.A(_3495_),
    .X(_3496_));
 sky130_fd_sc_hd__clkbuf_4 _3959_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_3497_));
 sky130_fd_sc_hd__nand2_1 _3960_ (.A(_3496_),
    .B(_3497_),
    .Y(_3498_));
 sky130_fd_sc_hd__o221a_1 _3961_ (.A1(_3488_),
    .A2(_3490_),
    .B1(_3491_),
    .B2(_3493_),
    .C1(_3498_),
    .X(_3499_));
 sky130_fd_sc_hd__inv_2 _3962_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_3500_));
 sky130_fd_sc_hd__nand2_2 _3963_ (.A(_3267_),
    .B(_3470_),
    .Y(_3501_));
 sky130_fd_sc_hd__buf_2 _3964_ (.A(_3501_),
    .X(_3502_));
 sky130_fd_sc_hd__inv_2 _3965_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .Y(_3503_));
 sky130_fd_sc_hd__nand2_2 _3966_ (.A(_3260_),
    .B(_3470_),
    .Y(_3504_));
 sky130_fd_sc_hd__buf_2 _3967_ (.A(_3504_),
    .X(_3505_));
 sky130_fd_sc_hd__o22ai_1 _3968_ (.A1(_3500_),
    .A2(_3502_),
    .B1(_3503_),
    .B2(_3505_),
    .Y(_3506_));
 sky130_fd_sc_hd__and2_2 _3969_ (.A(_3251_),
    .B(_3470_),
    .X(_3507_));
 sky130_fd_sc_hd__clkbuf_4 _3970_ (.A(_3507_),
    .X(_3508_));
 sky130_fd_sc_hd__clkbuf_4 _3971_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .X(_3509_));
 sky130_fd_sc_hd__and2_2 _3972_ (.A(_3119_),
    .B(_3470_),
    .X(_3510_));
 sky130_fd_sc_hd__clkbuf_4 _3973_ (.A(_3510_),
    .X(_3511_));
 sky130_fd_sc_hd__buf_2 _3974_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .X(_3512_));
 sky130_fd_sc_hd__a22o_1 _3975_ (.A1(_3508_),
    .A2(_3509_),
    .B1(_3511_),
    .B2(_3512_),
    .X(_3513_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(_3506_),
    .B(_3513_),
    .Y(_3514_));
 sky130_fd_sc_hd__and2_1 _3977_ (.A(_3307_),
    .B(_3469_),
    .X(_3515_));
 sky130_fd_sc_hd__clkbuf_2 _3978_ (.A(_3515_),
    .X(_0322_));
 sky130_fd_sc_hd__buf_2 _3979_ (.A(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_4 _3980_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_1 _3981_ (.A(_0323_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__and2_1 _3982_ (.A(_3316_),
    .B(_3469_),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_2 _3983_ (.A(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_4 _3984_ (.A(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _3985_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _3986_ (.A(_0328_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__and2_1 _3987_ (.A(_3302_),
    .B(_3469_),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_2 _3988_ (.A(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_4 _3989_ (.A(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_4 _3990_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _3991_ (.A(_0333_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__and2_1 _3992_ (.A(_3312_),
    .B(_3469_),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_2 _3993_ (.A(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__buf_4 _3994_ (.A(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_4 _3995_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_0338_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__and4_1 _3997_ (.A(_0325_),
    .B(_0330_),
    .C(_0335_),
    .D(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__and4_1 _3998_ (.A(_3487_),
    .B(_3499_),
    .C(_3514_),
    .D(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__and4_1 _3999_ (.A(_3321_),
    .B(_3394_),
    .C(_3467_),
    .D(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__and3_2 _4000_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_4 _4001_ (.A(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__and2_1 _4002_ (.A(_3242_),
    .B(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_2 _4003_ (.A(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__buf_2 _4004_ (.A(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__inv_2 _4005_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_2 _4006_ (.A(_3234_),
    .B(_0345_),
    .Y(_0350_));
 sky130_fd_sc_hd__clkbuf_4 _4007_ (.A(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_1 _4008_ (.A(_0349_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__and2_1 _4009_ (.A(_3217_),
    .B(_0345_),
    .X(_0353_));
 sky130_fd_sc_hd__buf_2 _4010_ (.A(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _4011_ (.A(_3226_),
    .B(_0345_),
    .X(_0355_));
 sky130_fd_sc_hd__buf_2 _4012_ (.A(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _4013_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .B1(_0356_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_0357_));
 sky130_fd_sc_hd__a211oi_1 _4014_ (.A1(_3174_),
    .A2(_0348_),
    .B1(_0352_),
    .C1(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__and2_1 _4015_ (.A(_3289_),
    .B(_0344_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_2 _4016_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_2 _4017_ (.A(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _4018_ (.A(_3292_),
    .B(_0345_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_2 _4019_ (.A(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_4 _4020_ (.A(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__inv_2 _4021_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_2 _4022_ (.A(_3278_),
    .B(_0345_),
    .Y(_0366_));
 sky130_fd_sc_hd__clkbuf_4 _4023_ (.A(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _4024_ (.A(_3283_),
    .B(_0344_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_2 _4025_ (.A(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__buf_2 _4026_ (.A(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_1 _4027_ (.A(_0370_),
    .B(_3163_),
    .Y(_0371_));
 sky130_fd_sc_hd__o21ai_1 _4028_ (.A1(_0365_),
    .A2(_0367_),
    .B1(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a221oi_1 _4029_ (.A1(_3168_),
    .A2(_0361_),
    .B1(_3171_),
    .B2(_0364_),
    .C1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__and2_1 _4030_ (.A(_3251_),
    .B(_0344_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_2 _4031_ (.A(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__buf_2 _4032_ (.A(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _4033_ (.A(_3119_),
    .B(_0345_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_2 _4034_ (.A(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_4 _4035_ (.A(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__inv_2 _4036_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_0380_));
 sky130_fd_sc_hd__nand2_2 _4037_ (.A(_3267_),
    .B(_0345_),
    .Y(_0381_));
 sky130_fd_sc_hd__buf_2 _4038_ (.A(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__inv_2 _4039_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .Y(_0383_));
 sky130_fd_sc_hd__nand2_2 _4040_ (.A(_3260_),
    .B(_0345_),
    .Y(_0384_));
 sky130_fd_sc_hd__buf_2 _4041_ (.A(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__o22ai_1 _4042_ (.A1(_0380_),
    .A2(_0382_),
    .B1(_0383_),
    .B2(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a221oi_1 _4043_ (.A1(_3205_),
    .A2(_0376_),
    .B1(_3208_),
    .B2(_0379_),
    .C1(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__and2_1 _4044_ (.A(_3312_),
    .B(_0344_),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_2 _4045_ (.A(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__buf_2 _4046_ (.A(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__and2_1 _4047_ (.A(_3316_),
    .B(_0344_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_2 _4048_ (.A(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__buf_2 _4049_ (.A(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__inv_2 _4050_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_0394_));
 sky130_fd_sc_hd__nand2_2 _4051_ (.A(_3307_),
    .B(_0345_),
    .Y(_0395_));
 sky130_fd_sc_hd__buf_2 _4052_ (.A(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _4053_ (.A(_3302_),
    .B(_0344_),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_2 _4054_ (.A(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_2 _4055_ (.A(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _4056_ (.A(_0399_),
    .B(_3192_),
    .Y(_0400_));
 sky130_fd_sc_hd__o21ai_1 _4057_ (.A1(_0394_),
    .A2(_0396_),
    .B1(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__a221oi_1 _4058_ (.A1(_3186_),
    .A2(_0390_),
    .B1(_3189_),
    .B2(_0393_),
    .C1(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__and4_1 _4059_ (.A(_0358_),
    .B(_0373_),
    .C(_0387_),
    .D(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__inv_2 _4060_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_0404_));
 sky130_fd_sc_hd__or3_2 _4061_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .B(_3120_),
    .C(_3218_),
    .X(_0405_));
 sky130_fd_sc_hd__inv_2 _4062_ (.A(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__buf_2 _4063_ (.A(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_2 _4064_ (.A(_3119_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__buf_2 _4065_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _4066_ (.A(_3267_),
    .B(_0407_),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_2 _4067_ (.A(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__buf_2 _4068_ (.A(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_4 _4069_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_1 _4070_ (.A(_0412_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__and2_1 _4071_ (.A(_3251_),
    .B(_0407_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_2 _4072_ (.A(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__buf_2 _4073_ (.A(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_4 _4074_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(_0417_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_2 _4076_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _4077_ (.A(_3260_),
    .B(_0407_),
    .Y(_0421_));
 sky130_fd_sc_hd__clkbuf_2 _4078_ (.A(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__or2_1 _4079_ (.A(_0420_),
    .B(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__o2111a_1 _4080_ (.A1(_0404_),
    .A2(_0409_),
    .B1(_0414_),
    .C1(_0419_),
    .D1(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__inv_2 _4081_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_0425_));
 sky130_fd_sc_hd__nand2_2 _4082_ (.A(_3226_),
    .B(_0407_),
    .Y(_0426_));
 sky130_fd_sc_hd__clkbuf_4 _4083_ (.A(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__and2_1 _4084_ (.A(_3242_),
    .B(_0406_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_2 _4085_ (.A(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_4 _4086_ (.A(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _4087_ (.A(_0430_),
    .B(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_0431_));
 sky130_fd_sc_hd__and2_1 _4088_ (.A(_3217_),
    .B(_0407_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_2 _4089_ (.A(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_4 _4090_ (.A(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_2 _4091_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .X(_0435_));
 sky130_fd_sc_hd__nand2_1 _4092_ (.A(_0434_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_2 _4093_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _4094_ (.A(_3234_),
    .B(_0407_),
    .Y(_0438_));
 sky130_fd_sc_hd__buf_2 _4095_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or2_1 _4096_ (.A(_0437_),
    .B(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__o2111a_1 _4097_ (.A1(_0425_),
    .A2(_0427_),
    .B1(_0431_),
    .C1(_0436_),
    .D1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_4 _4098_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .X(_0442_));
 sky130_fd_sc_hd__and2_1 _4099_ (.A(_3278_),
    .B(_0407_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_2 _4100_ (.A(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_4 _4101_ (.A(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_2 _4102_ (.A(_0405_),
    .B(_3282_),
    .Y(_0446_));
 sky130_fd_sc_hd__clkbuf_4 _4103_ (.A(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_4 _4104_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .X(_0448_));
 sky130_fd_sc_hd__and2_1 _4105_ (.A(_3292_),
    .B(_0406_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_2 _4106_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_2 _4107_ (.A(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_4 _4108_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_1 _4109_ (.A(_0451_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__and2_1 _4110_ (.A(_3289_),
    .B(_0406_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_2 _4111_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__buf_2 _4112_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_4 _4113_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_1 _4114_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand2_1 _4115_ (.A(_0453_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__a221oi_1 _4116_ (.A1(_0442_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0448_),
    .C1(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _4117_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .X(_0461_));
 sky130_fd_sc_hd__and2_1 _4118_ (.A(_3302_),
    .B(_0407_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_2 _4119_ (.A(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__buf_2 _4120_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__buf_2 _4121_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .X(_0465_));
 sky130_fd_sc_hd__and2_1 _4122_ (.A(_3307_),
    .B(_0407_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_2 _4123_ (.A(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_4 _4124_ (.A(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__and2_1 _4125_ (.A(_3316_),
    .B(_0406_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_2 _4126_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__buf_2 _4127_ (.A(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(_0471_),
    .B(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_0472_));
 sky130_fd_sc_hd__and2_1 _4129_ (.A(_3312_),
    .B(_0406_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_2 _4130_ (.A(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__buf_2 _4131_ (.A(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _4132_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(_0472_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__a221oi_1 _4134_ (.A1(_0461_),
    .A2(_0464_),
    .B1(_0465_),
    .B2(_0468_),
    .C1(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__and4_1 _4135_ (.A(_0424_),
    .B(_0441_),
    .C(_0460_),
    .D(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_1 _4136_ (.A(_0403_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_2 _4137_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0481_));
 sky130_fd_sc_hd__or3_2 _4138_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .B(_3120_),
    .C(_3396_),
    .X(_0482_));
 sky130_fd_sc_hd__inv_2 _4139_ (.A(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__clkbuf_4 _4140_ (.A(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__nand2_2 _4141_ (.A(_3234_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__clkbuf_4 _4142_ (.A(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__and2_1 _4143_ (.A(_3242_),
    .B(_0483_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_2 _4144_ (.A(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__buf_2 _4145_ (.A(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_1 _4146_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0490_));
 sky130_fd_sc_hd__o21ai_1 _4147_ (.A1(_0481_),
    .A2(_0486_),
    .B1(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__and2_1 _4148_ (.A(_3278_),
    .B(_0483_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_2 _4149_ (.A(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__buf_2 _4150_ (.A(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__nor2_2 _4151_ (.A(_0482_),
    .B(_3282_),
    .Y(_0495_));
 sky130_fd_sc_hd__buf_2 _4152_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__and2_1 _4153_ (.A(_3292_),
    .B(_0483_),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_2 _4154_ (.A(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__buf_2 _4155_ (.A(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_1 _4156_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0500_));
 sky130_fd_sc_hd__and2_1 _4157_ (.A(_3289_),
    .B(_0483_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_2 _4158_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__buf_4 _4159_ (.A(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__nand2_1 _4160_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_1 _4161_ (.A(_0500_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__a221oi_1 _4162_ (.A1(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .A2(_0494_),
    .B1(_0496_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .C1(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__and2_1 _4163_ (.A(_3217_),
    .B(_0484_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_2 _4164_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__buf_2 _4165_ (.A(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__buf_2 _4166_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _4167_ (.A(_0509_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__and2_1 _4168_ (.A(_3226_),
    .B(_0483_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_2 _4169_ (.A(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__buf_2 _4170_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__buf_2 _4171_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _4172_ (.A(_0514_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__and4b_1 _4173_ (.A_N(_0491_),
    .B(_0506_),
    .C(_0511_),
    .D(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_4 _4174_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_0518_));
 sky130_fd_sc_hd__and2_1 _4175_ (.A(_3302_),
    .B(_0484_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_2 _4176_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_4 _4177_ (.A(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_4 _4178_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_0522_));
 sky130_fd_sc_hd__and2_1 _4179_ (.A(_3307_),
    .B(_0484_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_2 _4180_ (.A(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_4 _4181_ (.A(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__inv_2 _4182_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_2 _4183_ (.A(_3312_),
    .B(_0484_),
    .Y(_0527_));
 sky130_fd_sc_hd__buf_2 _4184_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2_2 _4186_ (.A(_3316_),
    .B(_0484_),
    .Y(_0530_));
 sky130_fd_sc_hd__buf_2 _4187_ (.A(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__o22ai_1 _4188_ (.A1(_0526_),
    .A2(_0528_),
    .B1(_0529_),
    .B2(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__a221oi_1 _4189_ (.A1(_0518_),
    .A2(_0521_),
    .B1(_0522_),
    .B2(_0525_),
    .C1(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__buf_2 _4190_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .X(_0534_));
 sky130_fd_sc_hd__and2_1 _4191_ (.A(_3251_),
    .B(_0484_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_2 _4192_ (.A(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_4 _4193_ (.A(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_2 _4194_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .X(_0538_));
 sky130_fd_sc_hd__and2_1 _4195_ (.A(_3119_),
    .B(_0484_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_2 _4196_ (.A(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__clkbuf_4 _4197_ (.A(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__inv_2 _4198_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_2 _4199_ (.A(_3267_),
    .B(_0484_),
    .Y(_0543_));
 sky130_fd_sc_hd__buf_2 _4200_ (.A(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__inv_2 _4201_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_2 _4202_ (.A(_3260_),
    .B(_0484_),
    .Y(_0546_));
 sky130_fd_sc_hd__buf_2 _4203_ (.A(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o22ai_1 _4204_ (.A1(_0542_),
    .A2(_0544_),
    .B1(_0545_),
    .B2(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a221oi_1 _4205_ (.A1(_0534_),
    .A2(_0537_),
    .B1(_0538_),
    .B2(_0541_),
    .C1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__and3_1 _4206_ (.A(_0517_),
    .B(_0533_),
    .C(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_4 _4207_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_0551_));
 sky130_fd_sc_hd__and3_2 _4208_ (.A(_3396_),
    .B(_3218_),
    .C(\egd_top.BitStream_buffer.pc[6] ),
    .X(_0552_));
 sky130_fd_sc_hd__buf_2 _4209_ (.A(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__and2_1 _4210_ (.A(_3217_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_2 _4211_ (.A(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _4212_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__clkbuf_4 _4213_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_0557_));
 sky130_fd_sc_hd__and2_1 _4214_ (.A(_3226_),
    .B(_0553_),
    .X(_0558_));
 sky130_fd_sc_hd__clkbuf_2 _4215_ (.A(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__buf_2 _4216_ (.A(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__and2_1 _4217_ (.A(_3234_),
    .B(_0552_),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_2 _4218_ (.A(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__buf_2 _4219_ (.A(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_4 _4220_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _4221_ (.A(_0563_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__and2_1 _4222_ (.A(_3242_),
    .B(_0552_),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_2 _4223_ (.A(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__buf_2 _4224_ (.A(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__clkbuf_4 _4225_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_1 _4226_ (.A(_0568_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_1 _4227_ (.A(_0565_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__a221oi_1 _4228_ (.A1(_0551_),
    .A2(_0556_),
    .B1(_0557_),
    .B2(_0560_),
    .C1(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__buf_2 _4229_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_0573_));
 sky130_fd_sc_hd__and2_1 _4230_ (.A(_3251_),
    .B(_0553_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_2 _4231_ (.A(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_4 _4232_ (.A(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_4 _4233_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_0577_));
 sky130_fd_sc_hd__and2_1 _4234_ (.A(_3119_),
    .B(_0553_),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_2 _4235_ (.A(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_4 _4236_ (.A(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__and2_1 _4237_ (.A(_3260_),
    .B(_0552_),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_2 _4238_ (.A(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__buf_2 _4239_ (.A(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_4 _4240_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_0584_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(_0583_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__and2_1 _4242_ (.A(_3267_),
    .B(_0552_),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_2 _4243_ (.A(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__buf_2 _4244_ (.A(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_4 _4245_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_0589_));
 sky130_fd_sc_hd__nand2_1 _4246_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _4247_ (.A(_0585_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__a221oi_1 _4248_ (.A1(_0573_),
    .A2(_0576_),
    .B1(_0577_),
    .B2(_0580_),
    .C1(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__buf_2 _4249_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .X(_0593_));
 sky130_fd_sc_hd__and2_1 _4250_ (.A(_3289_),
    .B(_0553_),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_2 _4251_ (.A(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__buf_2 _4252_ (.A(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_4 _4253_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .X(_0597_));
 sky130_fd_sc_hd__and2_1 _4254_ (.A(_3292_),
    .B(_0553_),
    .X(_0598_));
 sky130_fd_sc_hd__clkbuf_2 _4255_ (.A(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__buf_2 _4256_ (.A(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__inv_2 _4257_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2_2 _4258_ (.A(_3278_),
    .B(_0553_),
    .Y(_0602_));
 sky130_fd_sc_hd__buf_2 _4259_ (.A(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__and2_1 _4260_ (.A(_3283_),
    .B(_0552_),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_2 _4261_ (.A(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__buf_2 _4262_ (.A(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_4 _4263_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_1 _4264_ (.A(_0606_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__o21ai_1 _4265_ (.A1(_0601_),
    .A2(_0603_),
    .B1(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__a221oi_1 _4266_ (.A1(_0593_),
    .A2(_0596_),
    .B1(_0597_),
    .B2(_0600_),
    .C1(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__clkbuf_4 _4267_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_0611_));
 sky130_fd_sc_hd__and2_1 _4268_ (.A(_3302_),
    .B(_0552_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_2 _4269_ (.A(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__buf_2 _4270_ (.A(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_4 _4271_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_0615_));
 sky130_fd_sc_hd__and2_1 _4272_ (.A(_3307_),
    .B(_0553_),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_2 _4273_ (.A(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_2 _4274_ (.A(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__inv_2 _4275_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_0619_));
 sky130_fd_sc_hd__nand2_2 _4276_ (.A(_3312_),
    .B(_0553_),
    .Y(_0620_));
 sky130_fd_sc_hd__buf_2 _4277_ (.A(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__inv_2 _4278_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_2 _4279_ (.A(_3316_),
    .B(_0553_),
    .Y(_0623_));
 sky130_fd_sc_hd__buf_2 _4280_ (.A(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__o22ai_1 _4281_ (.A1(_0619_),
    .A2(_0621_),
    .B1(_0622_),
    .B2(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__a221oi_1 _4282_ (.A1(_0611_),
    .A2(_0614_),
    .B1(_0615_),
    .B2(_0618_),
    .C1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__and4_1 _4283_ (.A(_0572_),
    .B(_0592_),
    .C(_0610_),
    .D(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_0550_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__nor2_1 _4285_ (.A(_0480_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__o41a_2 _4286_ (.A1(\egd_top.BitStream_buffer.pc[2] ),
    .A2(\egd_top.BitStream_buffer.pc[3] ),
    .A3(\egd_top.BitStream_buffer.pc[1] ),
    .A4(_3115_),
    .B1(_3470_),
    .X(_0630_));
 sky130_fd_sc_hd__and4b_1 _4287_ (.A_N(_0630_),
    .B(_3120_),
    .C(_3396_),
    .D(_3218_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_2 _4288_ (.A(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__buf_2 _4289_ (.A(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_4 _4290_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _4291_ (.A(_0633_),
    .B(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand3_2 _4292_ (.A(_0343_),
    .B(_0629_),
    .C(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__nor2_1 _4293_ (.A(_3212_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__nor2_1 _4294_ (.A(_3211_),
    .B(_0637_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21ai_1 _4295_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B1(_3081_),
    .Y(_0638_));
 sky130_fd_sc_hd__clkbuf_4 _4296_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .X(_0639_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(_3237_),
    .B(_3213_),
    .Y(_0640_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_3245_),
    .B(_3238_),
    .Y(_0641_));
 sky130_fd_sc_hd__nand2_1 _4299_ (.A(_0640_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__a221oi_1 _4300_ (.A1(_3224_),
    .A2(_3223_),
    .B1(_0639_),
    .B2(_3229_),
    .C1(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _4301_ (.A(_3263_),
    .B(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _4303_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__a221oi_1 _4304_ (.A1(_3255_),
    .A2(_3254_),
    .B1(_3432_),
    .B2(_3258_),
    .C1(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__clkbuf_4 _4305_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .X(_0648_));
 sky130_fd_sc_hd__inv_2 _4306_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _4307_ (.A(_3295_),
    .B(_3246_),
    .Y(_0650_));
 sky130_fd_sc_hd__o21ai_1 _4308_ (.A1(_0649_),
    .A2(_3291_),
    .B1(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__a221oi_1 _4309_ (.A1(_3287_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_0648_),
    .C1(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _4310_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .Y(_0653_));
 sky130_fd_sc_hd__o22ai_1 _4311_ (.A1(_3315_),
    .A2(_3314_),
    .B1(_0653_),
    .B2(_3318_),
    .Y(_0654_));
 sky130_fd_sc_hd__a221oi_1 _4312_ (.A1(_3306_),
    .A2(_3305_),
    .B1(_3271_),
    .B2(_3310_),
    .C1(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__and4_1 _4313_ (.A(_0643_),
    .B(_0647_),
    .C(_0652_),
    .D(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__buf_2 _4314_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .X(_0657_));
 sky130_fd_sc_hd__nand2_1 _4315_ (.A(_3335_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__o21ai_1 _4316_ (.A1(_0601_),
    .A2(_3332_),
    .B1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__a221oi_1 _4317_ (.A1(_3327_),
    .A2(_3326_),
    .B1(_3336_),
    .B2(_3330_),
    .C1(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _4318_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0661_));
 sky130_fd_sc_hd__buf_2 _4319_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(_3353_),
    .B(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__o21ai_1 _4321_ (.A1(_0661_),
    .A2(_3350_),
    .B1(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__a221oi_1 _4322_ (.A1(_3344_),
    .A2(_3343_),
    .B1(_3354_),
    .B2(_3347_),
    .C1(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__inv_2 _4323_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_0666_));
 sky130_fd_sc_hd__nand2_1 _4324_ (.A(_3371_),
    .B(_3358_),
    .Y(_0667_));
 sky130_fd_sc_hd__o21ai_1 _4325_ (.A1(_0666_),
    .A2(_3368_),
    .B1(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__a221oi_1 _4326_ (.A1(_3362_),
    .A2(_3361_),
    .B1(_3340_),
    .B2(_3365_),
    .C1(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _4327_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _4328_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _4329_ (.A(_0670_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__a221oi_1 _4330_ (.A1(_3380_),
    .A2(_3379_),
    .B1(_3322_),
    .B2(_3383_),
    .C1(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__and4_1 _4331_ (.A(_0660_),
    .B(_0665_),
    .C(_0669_),
    .D(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__buf_2 _4332_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_0675_));
 sky130_fd_sc_hd__inv_2 _4333_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .Y(_0676_));
 sky130_fd_sc_hd__o22ai_1 _4334_ (.A1(_3409_),
    .A2(_3408_),
    .B1(_0676_),
    .B2(_3411_),
    .Y(_0677_));
 sky130_fd_sc_hd__a221oi_1 _4335_ (.A1(_3402_),
    .A2(_3401_),
    .B1(_0675_),
    .B2(_3405_),
    .C1(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__buf_2 _4336_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_0679_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_3427_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__o21ai_1 _4338_ (.A1(_3366_),
    .A2(_3424_),
    .B1(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__a221oi_1 _4339_ (.A1(_3418_),
    .A2(_3417_),
    .B1(_3428_),
    .B2(_3421_),
    .C1(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__buf_2 _4340_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_0683_));
 sky130_fd_sc_hd__inv_2 _4341_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _4342_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_0685_));
 sky130_fd_sc_hd__o21ai_1 _4343_ (.A1(_0684_),
    .A2(_3442_),
    .B1(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__a221oi_1 _4344_ (.A1(_3439_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_0683_),
    .C1(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _4345_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2_1 _4346_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _4347_ (.A(_0688_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__a221oi_1 _4348_ (.A1(_3453_),
    .A2(_3452_),
    .B1(_3414_),
    .B2(_3456_),
    .C1(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__and4_1 _4349_ (.A(_0678_),
    .B(_0682_),
    .C(_0687_),
    .D(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__inv_2 _4350_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .Y(_0693_));
 sky130_fd_sc_hd__nand2_1 _4351_ (.A(_3475_),
    .B(_3482_),
    .Y(_0694_));
 sky130_fd_sc_hd__clkbuf_4 _4352_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_1 _4353_ (.A(_3480_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__inv_2 _4354_ (.A(_0339_),
    .Y(_0697_));
 sky130_fd_sc_hd__or2_1 _4355_ (.A(_0697_),
    .B(_3485_),
    .X(_0698_));
 sky130_fd_sc_hd__o2111a_1 _4356_ (.A1(_0693_),
    .A2(_3472_),
    .B1(_0694_),
    .C1(_0696_),
    .D1(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__inv_2 _4357_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .Y(_0700_));
 sky130_fd_sc_hd__clkbuf_4 _4358_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_1 _4359_ (.A(_3496_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__o221a_1 _4360_ (.A1(_0700_),
    .A2(_3490_),
    .B1(_3488_),
    .B2(_3493_),
    .C1(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__inv_2 _4361_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .Y(_0704_));
 sky130_fd_sc_hd__o22ai_1 _4362_ (.A1(_3503_),
    .A2(_3502_),
    .B1(_0704_),
    .B2(_3505_),
    .Y(_0705_));
 sky130_fd_sc_hd__a22o_1 _4363_ (.A1(_3508_),
    .A2(_3512_),
    .B1(_3511_),
    .B2(_3275_),
    .X(_0706_));
 sky130_fd_sc_hd__nor2_1 _4364_ (.A(_0705_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__clkbuf_4 _4365_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .X(_0708_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(_0323_),
    .B(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _4367_ (.A(_0328_),
    .B(_0334_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _4368_ (.A(_0333_),
    .B(_0324_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _4369_ (.A(_0338_),
    .B(_0329_),
    .Y(_0712_));
 sky130_fd_sc_hd__and4_1 _4370_ (.A(_0709_),
    .B(_0710_),
    .C(_0711_),
    .D(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__and4_1 _4371_ (.A(_0699_),
    .B(_0703_),
    .C(_0707_),
    .D(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__and4_1 _4372_ (.A(_0656_),
    .B(_0674_),
    .C(_0692_),
    .D(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__inv_2 _4373_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_0716_));
 sky130_fd_sc_hd__nor2_1 _4374_ (.A(_0716_),
    .B(_0351_),
    .Y(_0717_));
 sky130_fd_sc_hd__a22o_1 _4375_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .B1(_0356_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_0718_));
 sky130_fd_sc_hd__a211oi_1 _4376_ (.A1(_3177_),
    .A2(_0348_),
    .B1(_0717_),
    .C1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__inv_2 _4377_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_0720_));
 sky130_fd_sc_hd__nand2_1 _4378_ (.A(_0370_),
    .B(_3168_),
    .Y(_0721_));
 sky130_fd_sc_hd__o21ai_1 _4379_ (.A1(_0720_),
    .A2(_0367_),
    .B1(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__a221oi_1 _4380_ (.A1(_3171_),
    .A2(_0361_),
    .B1(_3174_),
    .B2(_0364_),
    .C1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__inv_2 _4381_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .Y(_0724_));
 sky130_fd_sc_hd__o22ai_1 _4382_ (.A1(_0383_),
    .A2(_0382_),
    .B1(_0724_),
    .B2(_0385_),
    .Y(_0725_));
 sky130_fd_sc_hd__a221oi_1 _4383_ (.A1(_3208_),
    .A2(_0376_),
    .B1(_0634_),
    .B2(_0379_),
    .C1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_1 _4384_ (.A(_0399_),
    .B(_3195_),
    .Y(_0727_));
 sky130_fd_sc_hd__o21ai_1 _4385_ (.A1(_0380_),
    .A2(_0396_),
    .B1(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__a221oi_1 _4386_ (.A1(_3189_),
    .A2(_0390_),
    .B1(_3192_),
    .B2(_0393_),
    .C1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__and4_1 _4387_ (.A(_0719_),
    .B(_0723_),
    .C(_0726_),
    .D(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__clkbuf_4 _4388_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .X(_0731_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(_0412_),
    .B(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__clkbuf_4 _4390_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .X(_0733_));
 sky130_fd_sc_hd__nand2_1 _4391_ (.A(_0417_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__inv_2 _4392_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_0735_));
 sky130_fd_sc_hd__or2_1 _4393_ (.A(_0735_),
    .B(_0422_),
    .X(_0736_));
 sky130_fd_sc_hd__o2111a_1 _4394_ (.A1(_0365_),
    .A2(_0409_),
    .B1(_0732_),
    .C1(_0734_),
    .D1(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__inv_2 _4395_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_0738_));
 sky130_fd_sc_hd__clkbuf_4 _4396_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_0739_));
 sky130_fd_sc_hd__nand2_1 _4397_ (.A(_0430_),
    .B(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__clkbuf_4 _4398_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_0741_));
 sky130_fd_sc_hd__nand2_1 _4399_ (.A(_0434_),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__inv_2 _4400_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_0743_));
 sky130_fd_sc_hd__or2_1 _4401_ (.A(_0743_),
    .B(_0439_),
    .X(_0744_));
 sky130_fd_sc_hd__o2111a_1 _4402_ (.A1(_0738_),
    .A2(_0427_),
    .B1(_0740_),
    .C1(_0742_),
    .D1(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_4 _4403_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_0746_));
 sky130_fd_sc_hd__nand2_1 _4404_ (.A(_0451_),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(_0456_),
    .B(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_0747_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__a221oi_1 _4407_ (.A1(_0448_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0457_),
    .C1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(_0471_),
    .B(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _4409_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _4410_ (.A(_0751_),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__a221oi_1 _4411_ (.A1(_0465_),
    .A2(_0464_),
    .B1(_0413_),
    .B2(_0468_),
    .C1(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__and4_1 _4412_ (.A(_0737_),
    .B(_0745_),
    .C(_0750_),
    .D(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__nand2_1 _4413_ (.A(_0730_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__inv_2 _4414_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2_1 _4415_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0758_));
 sky130_fd_sc_hd__o21ai_1 _4416_ (.A1(_0757_),
    .A2(_0486_),
    .B1(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__nand2_1 _4417_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _4418_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0761_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_0760_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__a221oi_1 _4420_ (.A1(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .A2(_0494_),
    .B1(_0496_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .C1(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_1 _4421_ (.A(_0509_),
    .B(_0515_),
    .Y(_0764_));
 sky130_fd_sc_hd__buf_2 _4422_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_0765_));
 sky130_fd_sc_hd__nand2_1 _4423_ (.A(_0514_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__and4b_1 _4424_ (.A_N(_0759_),
    .B(_0763_),
    .C(_0764_),
    .D(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__buf_2 _4425_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_0768_));
 sky130_fd_sc_hd__inv_2 _4426_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_0769_));
 sky130_fd_sc_hd__o22ai_1 _4427_ (.A1(_0529_),
    .A2(_0528_),
    .B1(_0769_),
    .B2(_0531_),
    .Y(_0770_));
 sky130_fd_sc_hd__a221oi_1 _4428_ (.A1(_0522_),
    .A2(_0521_),
    .B1(_0768_),
    .B2(_0525_),
    .C1(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__inv_2 _4429_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_0772_));
 sky130_fd_sc_hd__o22ai_1 _4430_ (.A1(_0545_),
    .A2(_0544_),
    .B1(_0772_),
    .B2(_0547_),
    .Y(_0773_));
 sky130_fd_sc_hd__a221oi_1 _4431_ (.A1(_0538_),
    .A2(_0537_),
    .B1(_0442_),
    .B2(_0541_),
    .C1(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__and3_1 _4432_ (.A(_0767_),
    .B(_0771_),
    .C(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__clkbuf_4 _4433_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_0776_));
 sky130_fd_sc_hd__nand2_1 _4434_ (.A(_0563_),
    .B(_0551_),
    .Y(_0777_));
 sky130_fd_sc_hd__nand2_1 _4435_ (.A(_0568_),
    .B(_0564_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand2_1 _4436_ (.A(_0777_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__a221oi_1 _4437_ (.A1(_0557_),
    .A2(_0556_),
    .B1(_0776_),
    .B2(_0560_),
    .C1(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__clkbuf_4 _4438_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _4439_ (.A(_0583_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_0782_));
 sky130_fd_sc_hd__nand2_1 _4440_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_0783_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(_0782_),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__a221oi_2 _4442_ (.A1(_0577_),
    .A2(_0576_),
    .B1(_0781_),
    .B2(_0580_),
    .C1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__inv_2 _4443_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _4444_ (.A(_0606_),
    .B(_0593_),
    .Y(_0787_));
 sky130_fd_sc_hd__o21ai_1 _4445_ (.A1(_0786_),
    .A2(_0603_),
    .B1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__a221oi_1 _4446_ (.A1(_0597_),
    .A2(_0596_),
    .B1(_0569_),
    .B2(_0600_),
    .C1(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _4447_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_0790_));
 sky130_fd_sc_hd__o22ai_1 _4448_ (.A1(_0622_),
    .A2(_0621_),
    .B1(_0790_),
    .B2(_0624_),
    .Y(_0791_));
 sky130_fd_sc_hd__a221oi_1 _4449_ (.A1(_0615_),
    .A2(_0614_),
    .B1(_0589_),
    .B2(_0618_),
    .C1(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__and4_1 _4450_ (.A(_0780_),
    .B(_0785_),
    .C(_0789_),
    .D(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _4451_ (.A(_0775_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__nor2_1 _4452_ (.A(_0756_),
    .B(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__clkbuf_4 _4453_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0796_));
 sky130_fd_sc_hd__nand2_1 _4454_ (.A(_0633_),
    .B(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__nand3_2 _4455_ (.A(_0715_),
    .B(_0795_),
    .C(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__nor2_1 _4456_ (.A(_3212_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__nor2_1 _4457_ (.A(_0638_),
    .B(_0799_),
    .Y(_0296_));
 sky130_fd_sc_hd__o21ai_1 _4458_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B1(_3081_),
    .Y(_0800_));
 sky130_fd_sc_hd__clkbuf_4 _4459_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .X(_0801_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_3237_),
    .B(_3224_),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_3245_),
    .B(_3213_),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(_0802_),
    .B(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__a221oi_1 _4463_ (.A1(_0639_),
    .A2(_3223_),
    .B1(_0801_),
    .B2(_3229_),
    .C1(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__nand2_1 _4464_ (.A(_3263_),
    .B(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2_1 _4465_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .Y(_0807_));
 sky130_fd_sc_hd__nand2_1 _4466_ (.A(_0806_),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__a221oi_1 _4467_ (.A1(_3432_),
    .A2(_3254_),
    .B1(_3439_),
    .B2(_3258_),
    .C1(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__inv_2 _4468_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _4469_ (.A(_3295_),
    .B(_3238_),
    .Y(_0811_));
 sky130_fd_sc_hd__o21ai_1 _4470_ (.A1(_0810_),
    .A2(_3291_),
    .B1(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__a221oi_2 _4471_ (.A1(_0648_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_3296_),
    .C1(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__inv_2 _4472_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .Y(_0814_));
 sky130_fd_sc_hd__o22ai_1 _4473_ (.A1(_0653_),
    .A2(_3314_),
    .B1(_0814_),
    .B2(_3318_),
    .Y(_0815_));
 sky130_fd_sc_hd__a221oi_1 _4474_ (.A1(_3271_),
    .A2(_3305_),
    .B1(_3264_),
    .B2(_3310_),
    .C1(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__and4_1 _4475_ (.A(_0805_),
    .B(_0809_),
    .C(_0813_),
    .D(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__buf_2 _4476_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .X(_0818_));
 sky130_fd_sc_hd__nand2_1 _4477_ (.A(_3335_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__o21ai_1 _4478_ (.A1(_0786_),
    .A2(_3332_),
    .B1(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a221oi_1 _4479_ (.A1(_3336_),
    .A2(_3326_),
    .B1(_0657_),
    .B2(_3330_),
    .C1(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _4480_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0822_));
 sky130_fd_sc_hd__clkbuf_4 _4481_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_3353_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__o21ai_1 _4483_ (.A1(_0822_),
    .A2(_3350_),
    .B1(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__a221oi_1 _4484_ (.A1(_3354_),
    .A2(_3343_),
    .B1(_0662_),
    .B2(_3347_),
    .C1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_2 _4485_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_0827_));
 sky130_fd_sc_hd__nand2_1 _4486_ (.A(_3371_),
    .B(_3362_),
    .Y(_0828_));
 sky130_fd_sc_hd__o21ai_1 _4487_ (.A1(_0827_),
    .A2(_3368_),
    .B1(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__a221oi_1 _4488_ (.A1(_3340_),
    .A2(_3361_),
    .B1(_3344_),
    .B2(_3365_),
    .C1(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand2_1 _4489_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .Y(_0831_));
 sky130_fd_sc_hd__nand2_1 _4490_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_1 _4491_ (.A(_0831_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__a221oi_2 _4492_ (.A1(_3322_),
    .A2(_3379_),
    .B1(_3327_),
    .B2(_3383_),
    .C1(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__and4_1 _4493_ (.A(_0821_),
    .B(_0826_),
    .C(_0830_),
    .D(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__buf_2 _4494_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0836_));
 sky130_fd_sc_hd__inv_2 _4495_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_0837_));
 sky130_fd_sc_hd__o22ai_1 _4496_ (.A1(_0676_),
    .A2(_3408_),
    .B1(_0837_),
    .B2(_3411_),
    .Y(_0838_));
 sky130_fd_sc_hd__a221oi_1 _4497_ (.A1(_0675_),
    .A2(_3401_),
    .B1(_0836_),
    .B2(_3405_),
    .C1(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__buf_2 _4498_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_3427_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__o21ai_1 _4500_ (.A1(_0666_),
    .A2(_3424_),
    .B1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__a221oi_1 _4501_ (.A1(_3428_),
    .A2(_3417_),
    .B1(_0679_),
    .B2(_3421_),
    .C1(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__clkbuf_4 _4502_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _4503_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .Y(_0845_));
 sky130_fd_sc_hd__o21ai_1 _4504_ (.A1(_3406_),
    .A2(_3442_),
    .B1(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__a221oi_1 _4505_ (.A1(_0683_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_0844_),
    .C1(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__nand2_1 _4506_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_0848_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_1 _4508_ (.A(_0848_),
    .B(_0849_),
    .Y(_0850_));
 sky130_fd_sc_hd__a221oi_1 _4509_ (.A1(_3414_),
    .A2(_3452_),
    .B1(_3418_),
    .B2(_3456_),
    .C1(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__and4_1 _4510_ (.A(_0839_),
    .B(_0843_),
    .C(_0847_),
    .D(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_3475_),
    .B(_0339_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_3480_),
    .B(_3476_),
    .Y(_0854_));
 sky130_fd_sc_hd__inv_2 _4513_ (.A(_0329_),
    .Y(_0855_));
 sky130_fd_sc_hd__or2_1 _4514_ (.A(_0855_),
    .B(_3485_),
    .X(_0856_));
 sky130_fd_sc_hd__o2111a_1 _4515_ (.A1(_3483_),
    .A2(_3472_),
    .B1(_0853_),
    .C1(_0854_),
    .D1(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__inv_2 _4516_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0858_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_3496_),
    .B(_0695_),
    .Y(_0859_));
 sky130_fd_sc_hd__o221a_1 _4518_ (.A1(_0858_),
    .A2(_3490_),
    .B1(_0700_),
    .B2(_3493_),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__inv_2 _4519_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .Y(_0861_));
 sky130_fd_sc_hd__o22ai_1 _4520_ (.A1(_0704_),
    .A2(_3502_),
    .B1(_0861_),
    .B2(_3505_),
    .Y(_0862_));
 sky130_fd_sc_hd__a22o_1 _4521_ (.A1(_3508_),
    .A2(_3275_),
    .B1(_3511_),
    .B2(_3287_),
    .X(_0863_));
 sky130_fd_sc_hd__nor2_1 _4522_ (.A(_0862_),
    .B(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__clkbuf_4 _4523_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .X(_0865_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_0323_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_0328_),
    .B(_0324_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(_0333_),
    .B(_0708_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand2_1 _4527_ (.A(_0338_),
    .B(_0334_),
    .Y(_0869_));
 sky130_fd_sc_hd__and4_1 _4528_ (.A(_0866_),
    .B(_0867_),
    .C(_0868_),
    .D(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__and4_1 _4529_ (.A(_0857_),
    .B(_0860_),
    .C(_0864_),
    .D(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__and4_1 _4530_ (.A(_0817_),
    .B(_0835_),
    .C(_0852_),
    .D(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__inv_2 _4531_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_1 _4532_ (.A(_0873_),
    .B(_0351_),
    .Y(_0874_));
 sky130_fd_sc_hd__a22o_1 _4533_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .B1(_0356_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_0875_));
 sky130_fd_sc_hd__a211oi_1 _4534_ (.A1(_3180_),
    .A2(_0348_),
    .B1(_0874_),
    .C1(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__inv_2 _4535_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_0877_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(_0370_),
    .B(_3171_),
    .Y(_0878_));
 sky130_fd_sc_hd__o21ai_1 _4537_ (.A1(_0877_),
    .A2(_0367_),
    .B1(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__a221oi_1 _4538_ (.A1(_3174_),
    .A2(_0361_),
    .B1(_3177_),
    .B2(_0364_),
    .C1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__inv_2 _4539_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .Y(_0881_));
 sky130_fd_sc_hd__o22ai_1 _4540_ (.A1(_0724_),
    .A2(_0382_),
    .B1(_0881_),
    .B2(_0385_),
    .Y(_0882_));
 sky130_fd_sc_hd__a221oi_1 _4541_ (.A1(_0634_),
    .A2(_0376_),
    .B1(_0796_),
    .B2(_0379_),
    .C1(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand2_1 _4542_ (.A(_0399_),
    .B(_3199_),
    .Y(_0884_));
 sky130_fd_sc_hd__o21ai_1 _4543_ (.A1(_0383_),
    .A2(_0396_),
    .B1(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__a221oi_1 _4544_ (.A1(_3192_),
    .A2(_0390_),
    .B1(_3195_),
    .B2(_0393_),
    .C1(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__and4_1 _4545_ (.A(_0876_),
    .B(_0880_),
    .C(_0883_),
    .D(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(_0412_),
    .B(_0418_),
    .Y(_0888_));
 sky130_fd_sc_hd__nand2_1 _4547_ (.A(_0417_),
    .B(_3152_),
    .Y(_0889_));
 sky130_fd_sc_hd__or2_1 _4548_ (.A(_0404_),
    .B(_0422_),
    .X(_0890_));
 sky130_fd_sc_hd__o2111a_1 _4549_ (.A1(_0720_),
    .A2(_0409_),
    .B1(_0888_),
    .C1(_0889_),
    .D1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__inv_2 _4550_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_1 _4551_ (.A(_0430_),
    .B(_0435_),
    .Y(_0893_));
 sky130_fd_sc_hd__clkbuf_4 _4552_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .X(_0894_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_0434_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2_1 _4554_ (.A(_0425_),
    .B(_0439_),
    .X(_0896_));
 sky130_fd_sc_hd__o2111a_1 _4555_ (.A1(_0892_),
    .A2(_0427_),
    .B1(_0893_),
    .C1(_0895_),
    .D1(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _4556_ (.A(_0451_),
    .B(_0739_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_0456_),
    .B(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_0898_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__a221oi_1 _4559_ (.A1(_0457_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0452_),
    .C1(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_0471_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_0902_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_0903_));
 sky130_fd_sc_hd__nand2_1 _4562_ (.A(_0902_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__a221oi_1 _4563_ (.A1(_0413_),
    .A2(_0464_),
    .B1(_0731_),
    .B2(_0468_),
    .C1(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__and4_1 _4564_ (.A(_0891_),
    .B(_0897_),
    .C(_0901_),
    .D(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__nand2_1 _4565_ (.A(_0887_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__inv_2 _4566_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_0908_));
 sky130_fd_sc_hd__nand2_1 _4567_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0909_));
 sky130_fd_sc_hd__o21ai_1 _4568_ (.A1(_0908_),
    .A2(_0486_),
    .B1(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2_1 _4569_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _4570_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0912_));
 sky130_fd_sc_hd__nand2_1 _4571_ (.A(_0911_),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__a221oi_1 _4572_ (.A1(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .A2(_0494_),
    .B1(_0496_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .C1(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand2_1 _4573_ (.A(_0509_),
    .B(_0765_),
    .Y(_0915_));
 sky130_fd_sc_hd__clkbuf_4 _4574_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_0514_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__and4b_1 _4576_ (.A_N(_0910_),
    .B(_0914_),
    .C(_0915_),
    .D(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__clkbuf_4 _4577_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0919_));
 sky130_fd_sc_hd__inv_2 _4578_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_0920_));
 sky130_fd_sc_hd__o22ai_1 _4579_ (.A1(_0769_),
    .A2(_0528_),
    .B1(_0920_),
    .B2(_0531_),
    .Y(_0921_));
 sky130_fd_sc_hd__a221oi_1 _4580_ (.A1(_0768_),
    .A2(_0521_),
    .B1(_0919_),
    .B2(_0525_),
    .C1(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__inv_2 _4581_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_0923_));
 sky130_fd_sc_hd__o22ai_1 _4582_ (.A1(_0772_),
    .A2(_0544_),
    .B1(_0923_),
    .B2(_0547_),
    .Y(_0924_));
 sky130_fd_sc_hd__a221oi_2 _4583_ (.A1(_0442_),
    .A2(_0537_),
    .B1(_0448_),
    .B2(_0541_),
    .C1(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__and3_1 _4584_ (.A(_0918_),
    .B(_0922_),
    .C(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_4 _4585_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_0927_));
 sky130_fd_sc_hd__nand2_1 _4586_ (.A(_0563_),
    .B(_0557_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand2_1 _4587_ (.A(_0568_),
    .B(_0551_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand2_1 _4588_ (.A(_0928_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__a221oi_1 _4589_ (.A1(_0776_),
    .A2(_0556_),
    .B1(_0927_),
    .B2(_0560_),
    .C1(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__clkbuf_4 _4590_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .X(_0932_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(_0583_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_1 _4592_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_0933_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__a221oi_1 _4594_ (.A1(_0781_),
    .A2(_0576_),
    .B1(_0932_),
    .B2(_0580_),
    .C1(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__inv_2 _4595_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _4596_ (.A(_0606_),
    .B(_0597_),
    .Y(_0938_));
 sky130_fd_sc_hd__o21ai_1 _4597_ (.A1(_0937_),
    .A2(_0603_),
    .B1(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__a221oi_1 _4598_ (.A1(_0569_),
    .A2(_0596_),
    .B1(_0564_),
    .B2(_0600_),
    .C1(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__inv_2 _4599_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_0941_));
 sky130_fd_sc_hd__o22ai_1 _4600_ (.A1(_0790_),
    .A2(_0621_),
    .B1(_0941_),
    .B2(_0624_),
    .Y(_0942_));
 sky130_fd_sc_hd__a221oi_1 _4601_ (.A1(_0589_),
    .A2(_0614_),
    .B1(_0584_),
    .B2(_0618_),
    .C1(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__and4_1 _4602_ (.A(_0931_),
    .B(_0936_),
    .C(_0940_),
    .D(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__nand2_1 _4603_ (.A(_0926_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__nor2_1 _4604_ (.A(_0907_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__clkbuf_4 _4605_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_0947_));
 sky130_fd_sc_hd__nand2_1 _4606_ (.A(_0633_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__nand3_1 _4607_ (.A(_0872_),
    .B(_0946_),
    .C(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__nor2_1 _4608_ (.A(_3212_),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_1 _4609_ (.A(_0800_),
    .B(_0950_),
    .Y(_0295_));
 sky130_fd_sc_hd__o21ai_1 _4610_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B1(_3081_),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_3237_),
    .B(_0639_),
    .Y(_0952_));
 sky130_fd_sc_hd__nand2_1 _4612_ (.A(_3245_),
    .B(_3224_),
    .Y(_0953_));
 sky130_fd_sc_hd__nand2_1 _4613_ (.A(_0952_),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__a221oi_1 _4614_ (.A1(_0801_),
    .A2(_3223_),
    .B1(_3300_),
    .B2(_3229_),
    .C1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _4615_ (.A(_3263_),
    .B(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_0956_));
 sky130_fd_sc_hd__nand2_1 _4616_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .Y(_0957_));
 sky130_fd_sc_hd__nand2_1 _4617_ (.A(_0956_),
    .B(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__a221oi_1 _4618_ (.A1(_3439_),
    .A2(_3254_),
    .B1(_0683_),
    .B2(_3258_),
    .C1(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_2 _4619_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .Y(_0960_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_3295_),
    .B(_3213_),
    .Y(_0961_));
 sky130_fd_sc_hd__o21ai_1 _4621_ (.A1(_0960_),
    .A2(_3291_),
    .B1(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__a221oi_1 _4622_ (.A1(_3296_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_3246_),
    .C1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__inv_2 _4623_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_0964_));
 sky130_fd_sc_hd__o22ai_1 _4624_ (.A1(_0814_),
    .A2(_3314_),
    .B1(_0964_),
    .B2(_3318_),
    .Y(_0965_));
 sky130_fd_sc_hd__a221oi_1 _4625_ (.A1(_3264_),
    .A2(_3305_),
    .B1(_3250_),
    .B2(_3310_),
    .C1(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__and4_1 _4626_ (.A(_0955_),
    .B(_0959_),
    .C(_0963_),
    .D(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__nand2_1 _4627_ (.A(_3335_),
    .B(_0607_),
    .Y(_0968_));
 sky130_fd_sc_hd__o21ai_1 _4628_ (.A1(_0937_),
    .A2(_3332_),
    .B1(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__a221oi_1 _4629_ (.A1(_0657_),
    .A2(_3326_),
    .B1(_0818_),
    .B2(_3330_),
    .C1(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__inv_2 _4630_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_0971_));
 sky130_fd_sc_hd__clkbuf_4 _4631_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .X(_0972_));
 sky130_fd_sc_hd__nand2_1 _4632_ (.A(_3353_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__o21ai_1 _4633_ (.A1(_0971_),
    .A2(_3350_),
    .B1(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__a221oi_1 _4634_ (.A1(_0662_),
    .A2(_3343_),
    .B1(_0823_),
    .B2(_3347_),
    .C1(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__inv_2 _4635_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_0976_));
 sky130_fd_sc_hd__nand2_1 _4636_ (.A(_3371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_0977_));
 sky130_fd_sc_hd__o21ai_1 _4637_ (.A1(_0976_),
    .A2(_3368_),
    .B1(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__a221oi_1 _4638_ (.A1(_3344_),
    .A2(_3361_),
    .B1(_3354_),
    .B2(_3365_),
    .C1(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__nand2_1 _4639_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .Y(_0980_));
 sky130_fd_sc_hd__nand2_1 _4640_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .Y(_0981_));
 sky130_fd_sc_hd__nand2_1 _4641_ (.A(_0980_),
    .B(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__a221oi_2 _4642_ (.A1(_3327_),
    .A2(_3379_),
    .B1(_3336_),
    .B2(_3383_),
    .C1(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__and4_1 _4643_ (.A(_0970_),
    .B(_0975_),
    .C(_0979_),
    .D(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__inv_2 _4644_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_0985_));
 sky130_fd_sc_hd__o22ai_1 _4645_ (.A1(_0837_),
    .A2(_3408_),
    .B1(_0985_),
    .B2(_3411_),
    .Y(_0986_));
 sky130_fd_sc_hd__a221oi_1 _4646_ (.A1(_0836_),
    .A2(_3401_),
    .B1(_3449_),
    .B2(_3405_),
    .C1(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand2_1 _4647_ (.A(_3427_),
    .B(_3372_),
    .Y(_0988_));
 sky130_fd_sc_hd__o21ai_1 _4648_ (.A1(_0827_),
    .A2(_3424_),
    .B1(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__a221oi_1 _4649_ (.A1(_0679_),
    .A2(_3417_),
    .B1(_0840_),
    .B2(_3421_),
    .C1(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__clkbuf_4 _4650_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_1 _4651_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .Y(_0992_));
 sky130_fd_sc_hd__o21ai_1 _4652_ (.A1(_3409_),
    .A2(_3442_),
    .B1(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__a221oi_1 _4653_ (.A1(_0844_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_0991_),
    .C1(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand2_1 _4654_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _4655_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_0996_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_0995_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__a221oi_1 _4657_ (.A1(_3418_),
    .A2(_3452_),
    .B1(_3428_),
    .B2(_3456_),
    .C1(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__and4_1 _4658_ (.A(_0987_),
    .B(_0990_),
    .C(_0994_),
    .D(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__nand2_1 _4659_ (.A(_3475_),
    .B(_0329_),
    .Y(_1000_));
 sky130_fd_sc_hd__nand2_1 _4660_ (.A(_3480_),
    .B(_3482_),
    .Y(_1001_));
 sky130_fd_sc_hd__inv_2 _4661_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_1002_));
 sky130_fd_sc_hd__or2_1 _4662_ (.A(_1002_),
    .B(_3485_),
    .X(_1003_));
 sky130_fd_sc_hd__o2111a_1 _4663_ (.A1(_0697_),
    .A2(_3472_),
    .B1(_1000_),
    .C1(_1001_),
    .D1(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__nand2_1 _4664_ (.A(_3496_),
    .B(_3476_),
    .Y(_1005_));
 sky130_fd_sc_hd__o221a_1 _4665_ (.A1(_3468_),
    .A2(_3490_),
    .B1(_0858_),
    .B2(_3493_),
    .C1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__inv_2 _4666_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1007_));
 sky130_fd_sc_hd__o22ai_1 _4667_ (.A1(_0861_),
    .A2(_3502_),
    .B1(_1007_),
    .B2(_3505_),
    .Y(_1008_));
 sky130_fd_sc_hd__a22o_1 _4668_ (.A1(_3508_),
    .A2(_3287_),
    .B1(_3511_),
    .B2(_0648_),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_1 _4669_ (.A(_1008_),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_0323_),
    .B(_3509_),
    .Y(_1011_));
 sky130_fd_sc_hd__nand2_1 _4671_ (.A(_0328_),
    .B(_0708_),
    .Y(_1012_));
 sky130_fd_sc_hd__nand2_1 _4672_ (.A(_0333_),
    .B(_0865_),
    .Y(_1013_));
 sky130_fd_sc_hd__nand2_1 _4673_ (.A(_0338_),
    .B(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1014_));
 sky130_fd_sc_hd__and4_1 _4674_ (.A(_1011_),
    .B(_1012_),
    .C(_1013_),
    .D(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__and4_1 _4675_ (.A(_1004_),
    .B(_1006_),
    .C(_1010_),
    .D(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__and4_1 _4676_ (.A(_0967_),
    .B(_0984_),
    .C(_0999_),
    .D(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__inv_2 _4677_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1018_));
 sky130_fd_sc_hd__nor2_1 _4678_ (.A(_1018_),
    .B(_0351_),
    .Y(_1019_));
 sky130_fd_sc_hd__a22o_1 _4679_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .B1(_0356_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_1020_));
 sky130_fd_sc_hd__a211oi_1 _4680_ (.A1(_3183_),
    .A2(_0348_),
    .B1(_1019_),
    .C1(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__inv_2 _4681_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_1022_));
 sky130_fd_sc_hd__nand2_1 _4682_ (.A(_0370_),
    .B(_3174_),
    .Y(_1023_));
 sky130_fd_sc_hd__o21ai_1 _4683_ (.A1(_1022_),
    .A2(_0367_),
    .B1(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__a221oi_1 _4684_ (.A1(_3177_),
    .A2(_0361_),
    .B1(_3180_),
    .B2(_0364_),
    .C1(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__inv_2 _4685_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1026_));
 sky130_fd_sc_hd__o22ai_1 _4686_ (.A1(_0881_),
    .A2(_0382_),
    .B1(_1026_),
    .B2(_0385_),
    .Y(_1027_));
 sky130_fd_sc_hd__a221oi_1 _4687_ (.A1(_0796_),
    .A2(_0376_),
    .B1(_0947_),
    .B2(_0379_),
    .C1(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(_0399_),
    .B(_3202_),
    .Y(_1029_));
 sky130_fd_sc_hd__o21ai_1 _4689_ (.A1(_0724_),
    .A2(_0396_),
    .B1(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__a221oi_1 _4690_ (.A1(_3195_),
    .A2(_0390_),
    .B1(_3199_),
    .B2(_0393_),
    .C1(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__and4_1 _4691_ (.A(_1021_),
    .B(_1025_),
    .C(_1028_),
    .D(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__nand2_1 _4692_ (.A(_0412_),
    .B(_0733_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _4693_ (.A(_0417_),
    .B(_3163_),
    .Y(_1034_));
 sky130_fd_sc_hd__or2_1 _4694_ (.A(_0365_),
    .B(_0422_),
    .X(_1035_));
 sky130_fd_sc_hd__o2111a_1 _4695_ (.A1(_0877_),
    .A2(_0409_),
    .B1(_1033_),
    .C1(_1034_),
    .D1(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__inv_2 _4696_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .Y(_1037_));
 sky130_fd_sc_hd__nand2_1 _4697_ (.A(_0430_),
    .B(_0741_),
    .Y(_1038_));
 sky130_fd_sc_hd__clkbuf_4 _4698_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .X(_1039_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(_0434_),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__or2_1 _4700_ (.A(_0738_),
    .B(_0439_),
    .X(_1041_));
 sky130_fd_sc_hd__o2111a_1 _4701_ (.A1(_1037_),
    .A2(_0427_),
    .B1(_1038_),
    .C1(_1040_),
    .D1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__nand2_1 _4702_ (.A(_0451_),
    .B(_0435_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _4703_ (.A(_0456_),
    .B(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_1044_));
 sky130_fd_sc_hd__nand2_1 _4704_ (.A(_1043_),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a221oi_1 _4705_ (.A1(_0452_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0746_),
    .C1(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__nand2_1 _4706_ (.A(_0471_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1047_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_1 _4708_ (.A(_1047_),
    .B(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__a221oi_1 _4709_ (.A1(_0731_),
    .A2(_0464_),
    .B1(_0418_),
    .B2(_0468_),
    .C1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__and4_1 _4710_ (.A(_1036_),
    .B(_1042_),
    .C(_1046_),
    .D(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__nand2_1 _4711_ (.A(_1032_),
    .B(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _4712_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1053_));
 sky130_fd_sc_hd__o21ai_1 _4713_ (.A1(_0526_),
    .A2(_0486_),
    .B1(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__clkbuf_4 _4714_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_1 _4715_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_1 _4716_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_1057_));
 sky130_fd_sc_hd__nand2_1 _4717_ (.A(_1056_),
    .B(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__a221oi_1 _4718_ (.A1(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_1055_),
    .C1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__nand2_1 _4719_ (.A(_0509_),
    .B(_0916_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand2_1 _4720_ (.A(_0514_),
    .B(_0518_),
    .Y(_1061_));
 sky130_fd_sc_hd__and4b_1 _4721_ (.A_N(_1054_),
    .B(_1059_),
    .C(_1060_),
    .D(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__o22ai_1 _4722_ (.A1(_0920_),
    .A2(_0528_),
    .B1(_0542_),
    .B2(_0531_),
    .Y(_1063_));
 sky130_fd_sc_hd__a221oi_1 _4723_ (.A1(_0919_),
    .A2(_0521_),
    .B1(_0534_),
    .B2(_0525_),
    .C1(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__inv_2 _4724_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_1065_));
 sky130_fd_sc_hd__o22ai_1 _4725_ (.A1(_0923_),
    .A2(_0544_),
    .B1(_1065_),
    .B2(_0547_),
    .Y(_1066_));
 sky130_fd_sc_hd__a221oi_1 _4726_ (.A1(_0448_),
    .A2(_0537_),
    .B1(_0457_),
    .B2(_0541_),
    .C1(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__and3_1 _4727_ (.A(_1062_),
    .B(_1064_),
    .C(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__nand2_1 _4728_ (.A(_0563_),
    .B(_0776_),
    .Y(_1069_));
 sky130_fd_sc_hd__nand2_1 _4729_ (.A(_0568_),
    .B(_0557_),
    .Y(_1070_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(_1069_),
    .B(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__a221oi_1 _4731_ (.A1(_0927_),
    .A2(_0556_),
    .B1(_0611_),
    .B2(_0560_),
    .C1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__buf_2 _4732_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .X(_1073_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_0583_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1074_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1075_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_1074_),
    .B(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__a221oi_2 _4736_ (.A1(_0932_),
    .A2(_0576_),
    .B1(_1073_),
    .B2(_0580_),
    .C1(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__inv_2 _4737_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_1078_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0606_),
    .B(_0569_),
    .Y(_1079_));
 sky130_fd_sc_hd__o21ai_1 _4739_ (.A1(_1078_),
    .A2(_0603_),
    .B1(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__a221oi_1 _4740_ (.A1(_0564_),
    .A2(_0596_),
    .B1(_0551_),
    .B2(_0600_),
    .C1(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__inv_2 _4741_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_1082_));
 sky130_fd_sc_hd__o22ai_1 _4742_ (.A1(_0941_),
    .A2(_0621_),
    .B1(_1082_),
    .B2(_0624_),
    .Y(_1083_));
 sky130_fd_sc_hd__a221oi_1 _4743_ (.A1(_0584_),
    .A2(_0614_),
    .B1(_0573_),
    .B2(_0618_),
    .C1(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__and4_1 _4744_ (.A(_1072_),
    .B(_1077_),
    .C(_1081_),
    .D(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__nand2_1 _4745_ (.A(_1068_),
    .B(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__nor2_1 _4746_ (.A(_1052_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_0633_),
    .B(_3497_),
    .Y(_1088_));
 sky130_fd_sc_hd__nand3_2 _4748_ (.A(_1017_),
    .B(_1087_),
    .C(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__nor2_1 _4749_ (.A(_3212_),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__nor2_1 _4750_ (.A(_0951_),
    .B(_1090_),
    .Y(_0294_));
 sky130_fd_sc_hd__o21ai_1 _4751_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(_3081_),
    .Y(_1091_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_3237_),
    .B(_0801_),
    .Y(_1092_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(_3245_),
    .B(_0639_),
    .Y(_1093_));
 sky130_fd_sc_hd__nand2_1 _4754_ (.A(_1092_),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__a221oi_1 _4755_ (.A1(_3300_),
    .A2(_3223_),
    .B1(_3306_),
    .B2(_3229_),
    .C1(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _4756_ (.A(_3263_),
    .B(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_1096_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_1097_));
 sky130_fd_sc_hd__nand2_1 _4758_ (.A(_1096_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__a221oi_1 _4759_ (.A1(_0683_),
    .A2(_3254_),
    .B1(_0844_),
    .B2(_3258_),
    .C1(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__inv_2 _4760_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _4761_ (.A(_3295_),
    .B(_3224_),
    .Y(_1101_));
 sky130_fd_sc_hd__o21ai_1 _4762_ (.A1(_1100_),
    .A2(_3291_),
    .B1(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__a221oi_1 _4763_ (.A1(_3246_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_3238_),
    .C1(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__inv_2 _4764_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_1104_));
 sky130_fd_sc_hd__o22ai_1 _4765_ (.A1(_0964_),
    .A2(_3314_),
    .B1(_1104_),
    .B2(_3318_),
    .Y(_1105_));
 sky130_fd_sc_hd__a221oi_1 _4766_ (.A1(_3250_),
    .A2(_3305_),
    .B1(_3255_),
    .B2(_3310_),
    .C1(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__and4_1 _4767_ (.A(_1095_),
    .B(_1099_),
    .C(_1103_),
    .D(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_3335_),
    .B(_0593_),
    .Y(_1108_));
 sky130_fd_sc_hd__o21ai_1 _4769_ (.A1(_1078_),
    .A2(_3332_),
    .B1(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__a221oi_1 _4770_ (.A1(_0818_),
    .A2(_3326_),
    .B1(_0607_),
    .B2(_3330_),
    .C1(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__inv_2 _4771_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_1 _4772_ (.A(_3353_),
    .B(_3376_),
    .Y(_1112_));
 sky130_fd_sc_hd__o21ai_1 _4773_ (.A1(_1111_),
    .A2(_3350_),
    .B1(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__a221oi_1 _4774_ (.A1(_0823_),
    .A2(_3343_),
    .B1(_0972_),
    .B2(_3347_),
    .C1(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__inv_2 _4775_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1115_));
 sky130_fd_sc_hd__nand2_1 _4776_ (.A(_3371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1116_));
 sky130_fd_sc_hd__o21ai_1 _4777_ (.A1(_1115_),
    .A2(_3368_),
    .B1(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__a221oi_1 _4778_ (.A1(_3354_),
    .A2(_3361_),
    .B1(_0662_),
    .B2(_3365_),
    .C1(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .Y(_1119_));
 sky130_fd_sc_hd__nand2_1 _4780_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .Y(_1120_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_1119_),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__a221oi_2 _4782_ (.A1(_3336_),
    .A2(_3379_),
    .B1(_0657_),
    .B2(_3383_),
    .C1(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__and4_1 _4783_ (.A(_1110_),
    .B(_1114_),
    .C(_1118_),
    .D(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__inv_2 _4784_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_1124_));
 sky130_fd_sc_hd__o22ai_1 _4785_ (.A1(_0985_),
    .A2(_3408_),
    .B1(_1124_),
    .B2(_3411_),
    .Y(_1125_));
 sky130_fd_sc_hd__a221oi_1 _4786_ (.A1(_3449_),
    .A2(_3401_),
    .B1(_3453_),
    .B2(_3405_),
    .C1(_1125_),
    .Y(_1126_));
 sky130_fd_sc_hd__nand2_1 _4787_ (.A(_3427_),
    .B(_3358_),
    .Y(_1127_));
 sky130_fd_sc_hd__o21ai_1 _4788_ (.A1(_0976_),
    .A2(_3424_),
    .B1(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__a221oi_1 _4789_ (.A1(_0840_),
    .A2(_3417_),
    .B1(_3372_),
    .B2(_3421_),
    .C1(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__clkbuf_4 _4790_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_1130_));
 sky130_fd_sc_hd__nand2_1 _4791_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_1131_));
 sky130_fd_sc_hd__o21ai_1 _4792_ (.A1(_0676_),
    .A2(_3442_),
    .B1(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__a221oi_1 _4793_ (.A1(_0991_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_1130_),
    .C1(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__nand2_1 _4794_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1134_));
 sky130_fd_sc_hd__nand2_1 _4795_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1135_));
 sky130_fd_sc_hd__nand2_1 _4796_ (.A(_1134_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__a221oi_1 _4797_ (.A1(_3428_),
    .A2(_3452_),
    .B1(_0679_),
    .B2(_3456_),
    .C1(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__and4_1 _4798_ (.A(_1126_),
    .B(_1129_),
    .C(_1133_),
    .D(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__nand2_1 _4799_ (.A(_3475_),
    .B(_0334_),
    .Y(_1139_));
 sky130_fd_sc_hd__nand2_1 _4800_ (.A(_3480_),
    .B(_0339_),
    .Y(_1140_));
 sky130_fd_sc_hd__inv_2 _4801_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_1141_));
 sky130_fd_sc_hd__or2_1 _4802_ (.A(_1141_),
    .B(_3485_),
    .X(_1142_));
 sky130_fd_sc_hd__o2111a_1 _4803_ (.A1(_0855_),
    .A2(_3472_),
    .B1(_1139_),
    .C1(_1140_),
    .D1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__nand2_1 _4804_ (.A(_3496_),
    .B(_3482_),
    .Y(_1144_));
 sky130_fd_sc_hd__o221a_1 _4805_ (.A1(_0693_),
    .A2(_3490_),
    .B1(_3468_),
    .B2(_3493_),
    .C1(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__inv_2 _4806_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_1146_));
 sky130_fd_sc_hd__o22ai_1 _4807_ (.A1(_1007_),
    .A2(_3502_),
    .B1(_1146_),
    .B2(_3505_),
    .Y(_1147_));
 sky130_fd_sc_hd__a22o_1 _4808_ (.A1(_3508_),
    .A2(_0648_),
    .B1(_3511_),
    .B2(_3296_),
    .X(_1148_));
 sky130_fd_sc_hd__nor2_1 _4809_ (.A(_1147_),
    .B(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _4810_ (.A(_0323_),
    .B(_3512_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_1 _4811_ (.A(_0328_),
    .B(_0865_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand2_1 _4812_ (.A(_0333_),
    .B(_3509_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _4813_ (.A(_0338_),
    .B(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_1153_));
 sky130_fd_sc_hd__and4_1 _4814_ (.A(_1150_),
    .B(_1151_),
    .C(_1152_),
    .D(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__and4_1 _4815_ (.A(_1143_),
    .B(_1145_),
    .C(_1149_),
    .D(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__and4_1 _4816_ (.A(_1107_),
    .B(_1123_),
    .C(_1138_),
    .D(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__inv_2 _4817_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1157_));
 sky130_fd_sc_hd__nor2_1 _4818_ (.A(_1157_),
    .B(_0351_),
    .Y(_1158_));
 sky130_fd_sc_hd__a22o_1 _4819_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .B1(_0356_),
    .B2(_3195_),
    .X(_1159_));
 sky130_fd_sc_hd__a211oi_1 _4820_ (.A1(_3186_),
    .A2(_0348_),
    .B1(_1158_),
    .C1(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__inv_2 _4821_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _4822_ (.A(_0370_),
    .B(_3177_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21ai_1 _4823_ (.A1(_1161_),
    .A2(_0367_),
    .B1(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__a221oi_1 _4824_ (.A1(_3180_),
    .A2(_0361_),
    .B1(_3183_),
    .B2(_0364_),
    .C1(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__o22ai_1 _4825_ (.A1(_1026_),
    .A2(_0382_),
    .B1(_3491_),
    .B2(_0385_),
    .Y(_1165_));
 sky130_fd_sc_hd__a221oi_2 _4826_ (.A1(_0947_),
    .A2(_0376_),
    .B1(_3497_),
    .B2(_0379_),
    .C1(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _4827_ (.A(_0399_),
    .B(_3205_),
    .Y(_1167_));
 sky130_fd_sc_hd__o21ai_1 _4828_ (.A1(_0881_),
    .A2(_0396_),
    .B1(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__a221oi_1 _4829_ (.A1(_3199_),
    .A2(_0390_),
    .B1(_3202_),
    .B2(_0393_),
    .C1(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__and4_1 _4830_ (.A(_1160_),
    .B(_1164_),
    .C(_1166_),
    .D(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nand2_1 _4831_ (.A(_0412_),
    .B(_3152_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_0417_),
    .B(_3168_),
    .Y(_1172_));
 sky130_fd_sc_hd__or2_1 _4833_ (.A(_0720_),
    .B(_0422_),
    .X(_1173_));
 sky130_fd_sc_hd__o2111a_1 _4834_ (.A1(_1022_),
    .A2(_0409_),
    .B1(_1171_),
    .C1(_1172_),
    .D1(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__inv_2 _4835_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _4836_ (.A(_0430_),
    .B(_0894_),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _4837_ (.A(_0434_),
    .B(_0461_),
    .Y(_1177_));
 sky130_fd_sc_hd__or2_1 _4838_ (.A(_0892_),
    .B(_0439_),
    .X(_1178_));
 sky130_fd_sc_hd__o2111a_1 _4839_ (.A1(_1175_),
    .A2(_0427_),
    .B1(_1176_),
    .C1(_1177_),
    .D1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__nand2_1 _4840_ (.A(_0451_),
    .B(_0741_),
    .Y(_1180_));
 sky130_fd_sc_hd__nand2_1 _4841_ (.A(_0456_),
    .B(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_1181_));
 sky130_fd_sc_hd__nand2_1 _4842_ (.A(_1180_),
    .B(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__a221oi_1 _4843_ (.A1(_0746_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0739_),
    .C1(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(_0471_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1184_));
 sky130_fd_sc_hd__nand2_1 _4845_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1185_));
 sky130_fd_sc_hd__nand2_1 _4846_ (.A(_1184_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__a221oi_1 _4847_ (.A1(_0418_),
    .A2(_0464_),
    .B1(_0733_),
    .B2(_0468_),
    .C1(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__and4_1 _4848_ (.A(_1174_),
    .B(_1179_),
    .C(_1183_),
    .D(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(_1170_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1190_));
 sky130_fd_sc_hd__o21ai_1 _4851_ (.A1(_0529_),
    .A2(_0486_),
    .B1(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__clkbuf_4 _4852_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_1192_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1193_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_1194_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_1193_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__a221oi_1 _4856_ (.A1(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_1192_),
    .C1(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(_0509_),
    .B(_0518_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_1 _4858_ (.A(_0514_),
    .B(_0522_),
    .Y(_1198_));
 sky130_fd_sc_hd__and4b_1 _4859_ (.A_N(_1191_),
    .B(_1196_),
    .C(_1197_),
    .D(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__o22ai_1 _4860_ (.A1(_0542_),
    .A2(_0528_),
    .B1(_0545_),
    .B2(_0531_),
    .Y(_1200_));
 sky130_fd_sc_hd__a221oi_1 _4861_ (.A1(_0534_),
    .A2(_0521_),
    .B1(_0538_),
    .B2(_0525_),
    .C1(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__inv_2 _4862_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_1202_));
 sky130_fd_sc_hd__o22ai_1 _4863_ (.A1(_1065_),
    .A2(_0544_),
    .B1(_1202_),
    .B2(_0547_),
    .Y(_1203_));
 sky130_fd_sc_hd__a221oi_1 _4864_ (.A1(_0457_),
    .A2(_0537_),
    .B1(_0452_),
    .B2(_0541_),
    .C1(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__and3_1 _4865_ (.A(_1199_),
    .B(_1201_),
    .C(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__nand2_1 _4866_ (.A(_0563_),
    .B(_0927_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(_0568_),
    .B(_0776_),
    .Y(_1207_));
 sky130_fd_sc_hd__nand2_1 _4868_ (.A(_1206_),
    .B(_1207_),
    .Y(_1208_));
 sky130_fd_sc_hd__a221oi_1 _4869_ (.A1(_0611_),
    .A2(_0556_),
    .B1(_0615_),
    .B2(_0560_),
    .C1(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__clkbuf_4 _4870_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .X(_1210_));
 sky130_fd_sc_hd__nand2_1 _4871_ (.A(_0583_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1211_));
 sky130_fd_sc_hd__nand2_1 _4872_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_1211_),
    .B(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__a221oi_1 _4874_ (.A1(_1073_),
    .A2(_0576_),
    .B1(_1210_),
    .B2(_0580_),
    .C1(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__inv_2 _4875_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_1 _4876_ (.A(_0606_),
    .B(_0564_),
    .Y(_1216_));
 sky130_fd_sc_hd__o21ai_1 _4877_ (.A1(_1215_),
    .A2(_0603_),
    .B1(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__a221oi_1 _4878_ (.A1(_0551_),
    .A2(_0596_),
    .B1(_0557_),
    .B2(_0600_),
    .C1(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__inv_2 _4879_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1219_));
 sky130_fd_sc_hd__o22ai_1 _4880_ (.A1(_1082_),
    .A2(_0621_),
    .B1(_1219_),
    .B2(_0624_),
    .Y(_1220_));
 sky130_fd_sc_hd__a221oi_1 _4881_ (.A1(_0573_),
    .A2(_0614_),
    .B1(_0577_),
    .B2(_0618_),
    .C1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__and4_1 _4882_ (.A(_1209_),
    .B(_1214_),
    .C(_1218_),
    .D(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__nand2_1 _4883_ (.A(_1205_),
    .B(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__nor2_1 _4884_ (.A(_1189_),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(_0633_),
    .B(_0701_),
    .Y(_1225_));
 sky130_fd_sc_hd__nand3_2 _4886_ (.A(_1156_),
    .B(_1224_),
    .C(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__nor2_1 _4887_ (.A(_3212_),
    .B(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__nor2_1 _4888_ (.A(_1091_),
    .B(_1227_),
    .Y(_0293_));
 sky130_fd_sc_hd__o21ai_1 _4889_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B1(_3081_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(_3237_),
    .B(_3300_),
    .Y(_1229_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_3245_),
    .B(_0801_),
    .Y(_1230_));
 sky130_fd_sc_hd__nand2_1 _4892_ (.A(_1229_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__a221oi_1 _4893_ (.A1(_3306_),
    .A2(_3223_),
    .B1(_3271_),
    .B2(_3229_),
    .C1(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2_1 _4894_ (.A(_3263_),
    .B(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_1233_));
 sky130_fd_sc_hd__nand2_1 _4895_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_1234_));
 sky130_fd_sc_hd__nand2_1 _4896_ (.A(_1233_),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__a221oi_1 _4897_ (.A1(_0844_),
    .A2(_3254_),
    .B1(_0991_),
    .B2(_3258_),
    .C1(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__inv_2 _4898_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _4899_ (.A(_3295_),
    .B(_0639_),
    .Y(_1238_));
 sky130_fd_sc_hd__o21ai_1 _4900_ (.A1(_1237_),
    .A2(_3291_),
    .B1(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__a221oi_1 _4901_ (.A1(_3238_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_3213_),
    .C1(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__inv_2 _4902_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .Y(_1241_));
 sky130_fd_sc_hd__o22ai_1 _4903_ (.A1(_1104_),
    .A2(_3314_),
    .B1(_1241_),
    .B2(_3318_),
    .Y(_1242_));
 sky130_fd_sc_hd__a221oi_1 _4904_ (.A1(_3255_),
    .A2(_3305_),
    .B1(_3432_),
    .B2(_3310_),
    .C1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__and4_1 _4905_ (.A(_1232_),
    .B(_1236_),
    .C(_1240_),
    .D(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(_3335_),
    .B(_0597_),
    .Y(_1245_));
 sky130_fd_sc_hd__o21ai_1 _4907_ (.A1(_1215_),
    .A2(_3332_),
    .B1(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a221oi_1 _4908_ (.A1(_0607_),
    .A2(_3326_),
    .B1(_0593_),
    .B2(_3330_),
    .C1(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__inv_2 _4909_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .Y(_1248_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(_3353_),
    .B(_3380_),
    .Y(_1249_));
 sky130_fd_sc_hd__o21ai_1 _4911_ (.A1(_1248_),
    .A2(_3350_),
    .B1(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__a221oi_1 _4912_ (.A1(_0972_),
    .A2(_3343_),
    .B1(_3376_),
    .B2(_3347_),
    .C1(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__inv_2 _4913_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_1 _4914_ (.A(_3371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1253_));
 sky130_fd_sc_hd__o21ai_1 _4915_ (.A1(_1252_),
    .A2(_3368_),
    .B1(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__a221oi_1 _4916_ (.A1(_0662_),
    .A2(_3361_),
    .B1(_0823_),
    .B2(_3365_),
    .C1(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__nand2_1 _4917_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _4918_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .Y(_1257_));
 sky130_fd_sc_hd__nand2_1 _4919_ (.A(_1256_),
    .B(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__a221oi_1 _4920_ (.A1(_0657_),
    .A2(_3379_),
    .B1(_0818_),
    .B2(_3383_),
    .C1(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__and4_1 _4921_ (.A(_1247_),
    .B(_1251_),
    .C(_1255_),
    .D(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__inv_2 _4922_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1261_));
 sky130_fd_sc_hd__o22ai_1 _4923_ (.A1(_1124_),
    .A2(_3408_),
    .B1(_1261_),
    .B2(_3411_),
    .Y(_1262_));
 sky130_fd_sc_hd__a221oi_1 _4924_ (.A1(_3453_),
    .A2(_3401_),
    .B1(_3414_),
    .B2(_3405_),
    .C1(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _4925_ (.A(_3427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_1264_));
 sky130_fd_sc_hd__o21ai_1 _4926_ (.A1(_1115_),
    .A2(_3424_),
    .B1(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__a221oi_1 _4927_ (.A1(_3372_),
    .A2(_3417_),
    .B1(_3358_),
    .B2(_3421_),
    .C1(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_1267_));
 sky130_fd_sc_hd__o21ai_1 _4929_ (.A1(_0837_),
    .A2(_3442_),
    .B1(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hd__a221oi_1 _4930_ (.A1(_1130_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_3395_),
    .C1(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__nand2_1 _4931_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1270_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1271_));
 sky130_fd_sc_hd__nand2_1 _4933_ (.A(_1270_),
    .B(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__a221oi_1 _4934_ (.A1(_0679_),
    .A2(_3452_),
    .B1(_0840_),
    .B2(_3456_),
    .C1(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__and4_1 _4935_ (.A(_1263_),
    .B(_1266_),
    .C(_1269_),
    .D(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(_3475_),
    .B(_0324_),
    .Y(_1275_));
 sky130_fd_sc_hd__nand2_1 _4937_ (.A(_3480_),
    .B(_0329_),
    .Y(_1276_));
 sky130_fd_sc_hd__or2_1 _4938_ (.A(_3500_),
    .B(_3485_),
    .X(_1277_));
 sky130_fd_sc_hd__o2111a_1 _4939_ (.A1(_1002_),
    .A2(_3472_),
    .B1(_1275_),
    .C1(_1276_),
    .D1(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_3496_),
    .B(_0339_),
    .Y(_1279_));
 sky130_fd_sc_hd__o221a_1 _4941_ (.A1(_3483_),
    .A2(_3490_),
    .B1(_0693_),
    .B2(_3493_),
    .C1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__o22ai_1 _4942_ (.A1(_1146_),
    .A2(_3502_),
    .B1(_3288_),
    .B2(_3505_),
    .Y(_1281_));
 sky130_fd_sc_hd__a22o_1 _4943_ (.A1(_3508_),
    .A2(_3296_),
    .B1(_3511_),
    .B2(_3246_),
    .X(_1282_));
 sky130_fd_sc_hd__nor2_1 _4944_ (.A(_1281_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__nand2_1 _4945_ (.A(_0323_),
    .B(_3275_),
    .Y(_1284_));
 sky130_fd_sc_hd__nand2_1 _4946_ (.A(_0328_),
    .B(_3509_),
    .Y(_1285_));
 sky130_fd_sc_hd__nand2_1 _4947_ (.A(_0333_),
    .B(_3512_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_1 _4948_ (.A(_0338_),
    .B(_0865_),
    .Y(_1287_));
 sky130_fd_sc_hd__and4_1 _4949_ (.A(_1284_),
    .B(_1285_),
    .C(_1286_),
    .D(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__and4_1 _4950_ (.A(_1278_),
    .B(_1280_),
    .C(_1283_),
    .D(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__and4_1 _4951_ (.A(_1244_),
    .B(_1260_),
    .C(_1274_),
    .D(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__inv_2 _4952_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1291_));
 sky130_fd_sc_hd__nor2_1 _4953_ (.A(_1291_),
    .B(_0351_),
    .Y(_1292_));
 sky130_fd_sc_hd__a22o_1 _4954_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .B1(_0356_),
    .B2(_3199_),
    .X(_1293_));
 sky130_fd_sc_hd__a211oi_1 _4955_ (.A1(_3189_),
    .A2(_0348_),
    .B1(_1292_),
    .C1(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__nand2_1 _4956_ (.A(_0370_),
    .B(_3180_),
    .Y(_1295_));
 sky130_fd_sc_hd__o21ai_1 _4957_ (.A1(_0349_),
    .A2(_0367_),
    .B1(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__a221oi_1 _4958_ (.A1(_3183_),
    .A2(_0361_),
    .B1(_3186_),
    .B2(_0364_),
    .C1(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__o22ai_1 _4959_ (.A1(_3491_),
    .A2(_0382_),
    .B1(_3488_),
    .B2(_0385_),
    .Y(_1298_));
 sky130_fd_sc_hd__a221oi_1 _4960_ (.A1(_3497_),
    .A2(_0376_),
    .B1(_0701_),
    .B2(_0379_),
    .C1(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _4961_ (.A(_0399_),
    .B(_3208_),
    .Y(_1300_));
 sky130_fd_sc_hd__o21ai_1 _4962_ (.A1(_1026_),
    .A2(_0396_),
    .B1(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__a221oi_1 _4963_ (.A1(_3202_),
    .A2(_0390_),
    .B1(_3205_),
    .B2(_0393_),
    .C1(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__and4_1 _4964_ (.A(_1294_),
    .B(_1297_),
    .C(_1299_),
    .D(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__nand2_1 _4965_ (.A(_0412_),
    .B(_3163_),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _4966_ (.A(_0417_),
    .B(_3171_),
    .Y(_1305_));
 sky130_fd_sc_hd__or2_1 _4967_ (.A(_0877_),
    .B(_0422_),
    .X(_1306_));
 sky130_fd_sc_hd__o2111a_1 _4968_ (.A1(_1161_),
    .A2(_0409_),
    .B1(_1304_),
    .C1(_1305_),
    .D1(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__inv_2 _4969_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1308_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_0430_),
    .B(_1039_),
    .Y(_1309_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_0434_),
    .B(_0465_),
    .Y(_1310_));
 sky130_fd_sc_hd__or2_1 _4972_ (.A(_1037_),
    .B(_0439_),
    .X(_1311_));
 sky130_fd_sc_hd__o2111a_1 _4973_ (.A1(_1308_),
    .A2(_0427_),
    .B1(_1309_),
    .C1(_1310_),
    .D1(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_0451_),
    .B(_0894_),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2_1 _4975_ (.A(_0456_),
    .B(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .Y(_1314_));
 sky130_fd_sc_hd__nand2_1 _4976_ (.A(_1313_),
    .B(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__a221oi_1 _4977_ (.A1(_0739_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0435_),
    .C1(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(_0471_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1317_));
 sky130_fd_sc_hd__nand2_1 _4979_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_1318_));
 sky130_fd_sc_hd__nand2_1 _4980_ (.A(_1317_),
    .B(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__a221oi_1 _4981_ (.A1(_0733_),
    .A2(_0464_),
    .B1(_3152_),
    .B2(_0468_),
    .C1(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__and4_1 _4982_ (.A(_1307_),
    .B(_1312_),
    .C(_1316_),
    .D(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__nand2_1 _4983_ (.A(_1303_),
    .B(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__nand2_1 _4984_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_1323_));
 sky130_fd_sc_hd__o21ai_1 _4985_ (.A1(_0769_),
    .A2(_0486_),
    .B1(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _4986_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _4987_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1326_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_1325_),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__a221oi_1 _4989_ (.A1(_1192_),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0510_),
    .C1(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2_1 _4990_ (.A(_0509_),
    .B(_0522_),
    .Y(_1329_));
 sky130_fd_sc_hd__nand2_1 _4991_ (.A(_0514_),
    .B(_0768_),
    .Y(_1330_));
 sky130_fd_sc_hd__and4b_1 _4992_ (.A_N(_1324_),
    .B(_1328_),
    .C(_1329_),
    .D(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__o22ai_1 _4993_ (.A1(_0545_),
    .A2(_0528_),
    .B1(_0772_),
    .B2(_0531_),
    .Y(_1332_));
 sky130_fd_sc_hd__a221oi_1 _4994_ (.A1(_0538_),
    .A2(_0521_),
    .B1(_0442_),
    .B2(_0525_),
    .C1(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__inv_2 _4995_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .Y(_1334_));
 sky130_fd_sc_hd__o22ai_1 _4996_ (.A1(_1202_),
    .A2(_0544_),
    .B1(_1334_),
    .B2(_0547_),
    .Y(_1335_));
 sky130_fd_sc_hd__a221oi_1 _4997_ (.A1(_0452_),
    .A2(_0537_),
    .B1(_0746_),
    .B2(_0541_),
    .C1(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hd__and3_1 _4998_ (.A(_1331_),
    .B(_1333_),
    .C(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__nand2_1 _4999_ (.A(_0563_),
    .B(_0611_),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _5000_ (.A(_0568_),
    .B(_0927_),
    .Y(_1339_));
 sky130_fd_sc_hd__nand2_1 _5001_ (.A(_1338_),
    .B(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__a221oi_1 _5002_ (.A1(_0615_),
    .A2(_0556_),
    .B1(_0589_),
    .B2(_0560_),
    .C1(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _5003_ (.A(_0583_),
    .B(_1073_),
    .Y(_1342_));
 sky130_fd_sc_hd__nand2_1 _5004_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1343_));
 sky130_fd_sc_hd__nand2_1 _5005_ (.A(_1342_),
    .B(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__a221oi_2 _5006_ (.A1(_1210_),
    .A2(_0576_),
    .B1(_1055_),
    .B2(_0580_),
    .C1(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__inv_2 _5007_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_1346_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1347_));
 sky130_fd_sc_hd__o21ai_1 _5009_ (.A1(_1346_),
    .A2(_0603_),
    .B1(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__a221oi_1 _5010_ (.A1(_0557_),
    .A2(_0596_),
    .B1(_0776_),
    .B2(_0600_),
    .C1(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__inv_2 _5011_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_1350_));
 sky130_fd_sc_hd__o22ai_1 _5012_ (.A1(_1219_),
    .A2(_0621_),
    .B1(_1350_),
    .B2(_0624_),
    .Y(_1351_));
 sky130_fd_sc_hd__a221oi_1 _5013_ (.A1(_0577_),
    .A2(_0614_),
    .B1(_0781_),
    .B2(_0618_),
    .C1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__and4_1 _5014_ (.A(_1341_),
    .B(_1345_),
    .C(_1349_),
    .D(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__nand2_1 _5015_ (.A(_1337_),
    .B(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__nor2_1 _5016_ (.A(_1322_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_1 _5017_ (.A(_0633_),
    .B(_0695_),
    .Y(_1356_));
 sky130_fd_sc_hd__nand3_2 _5018_ (.A(_1290_),
    .B(_1355_),
    .C(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__nor2_1 _5019_ (.A(_3212_),
    .B(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__nor2_1 _5020_ (.A(_1228_),
    .B(_1358_),
    .Y(_0292_));
 sky130_fd_sc_hd__o21ai_1 _5021_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B1(_3161_),
    .Y(_1359_));
 sky130_fd_sc_hd__nand2_1 _5022_ (.A(_3237_),
    .B(_3306_),
    .Y(_1360_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(_3245_),
    .B(_3300_),
    .Y(_1361_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(_1360_),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__a221oi_1 _5025_ (.A1(_3271_),
    .A2(_3223_),
    .B1(_3264_),
    .B2(_3229_),
    .C1(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_3263_),
    .B(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_1364_));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_1365_));
 sky130_fd_sc_hd__nand2_1 _5028_ (.A(_1364_),
    .B(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__a221oi_1 _5029_ (.A1(_0991_),
    .A2(_3254_),
    .B1(_1130_),
    .B2(_3258_),
    .C1(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_3295_),
    .B(_0801_),
    .Y(_1368_));
 sky130_fd_sc_hd__o21ai_1 _5031_ (.A1(_3311_),
    .A2(_3291_),
    .B1(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__a221oi_1 _5032_ (.A1(_3213_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_3224_),
    .C1(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__inv_2 _5033_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .Y(_1371_));
 sky130_fd_sc_hd__o22ai_1 _5034_ (.A1(_1241_),
    .A2(_3314_),
    .B1(_1371_),
    .B2(_3318_),
    .Y(_1372_));
 sky130_fd_sc_hd__a221oi_1 _5035_ (.A1(_3432_),
    .A2(_3305_),
    .B1(_3439_),
    .B2(_3310_),
    .C1(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__and4_1 _5036_ (.A(_1363_),
    .B(_1367_),
    .C(_1370_),
    .D(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__nand2_1 _5037_ (.A(_3335_),
    .B(_0569_),
    .Y(_1375_));
 sky130_fd_sc_hd__o21ai_1 _5038_ (.A1(_1346_),
    .A2(_3332_),
    .B1(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__a221oi_1 _5039_ (.A1(_0593_),
    .A2(_3326_),
    .B1(_0597_),
    .B2(_3330_),
    .C1(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__inv_2 _5040_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _5041_ (.A(_3353_),
    .B(_3322_),
    .Y(_1379_));
 sky130_fd_sc_hd__o21ai_1 _5042_ (.A1(_1378_),
    .A2(_3350_),
    .B1(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__a221oi_1 _5043_ (.A1(_3376_),
    .A2(_3343_),
    .B1(_3380_),
    .B2(_3347_),
    .C1(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__inv_2 _5044_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _5045_ (.A(_3371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1383_));
 sky130_fd_sc_hd__o21ai_1 _5046_ (.A1(_1382_),
    .A2(_3368_),
    .B1(_1383_),
    .Y(_1384_));
 sky130_fd_sc_hd__a221oi_1 _5047_ (.A1(_0823_),
    .A2(_3361_),
    .B1(_0972_),
    .B2(_3365_),
    .C1(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_1386_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_1387_));
 sky130_fd_sc_hd__nand2_1 _5050_ (.A(_1386_),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__a221oi_1 _5051_ (.A1(_0818_),
    .A2(_3379_),
    .B1(_0607_),
    .B2(_3383_),
    .C1(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__and4_1 _5052_ (.A(_1377_),
    .B(_1381_),
    .C(_1385_),
    .D(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__inv_2 _5053_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_1391_));
 sky130_fd_sc_hd__o22ai_1 _5054_ (.A1(_1261_),
    .A2(_3408_),
    .B1(_1391_),
    .B2(_3411_),
    .Y(_1392_));
 sky130_fd_sc_hd__a221oi_1 _5055_ (.A1(_3414_),
    .A2(_3401_),
    .B1(_3418_),
    .B2(_3405_),
    .C1(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2_1 _5056_ (.A(_3427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_1394_));
 sky130_fd_sc_hd__o21ai_1 _5057_ (.A1(_1252_),
    .A2(_3424_),
    .B1(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__a221oi_1 _5058_ (.A1(_3358_),
    .A2(_3417_),
    .B1(_3362_),
    .B2(_3421_),
    .C1(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__nand2_1 _5059_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .Y(_1397_));
 sky130_fd_sc_hd__o21ai_1 _5060_ (.A1(_0985_),
    .A2(_3442_),
    .B1(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__a221oi_1 _5061_ (.A1(_3395_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_3402_),
    .C1(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__nand2_1 _5062_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_1400_));
 sky130_fd_sc_hd__nand2_1 _5063_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1401_));
 sky130_fd_sc_hd__nand2_1 _5064_ (.A(_1400_),
    .B(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__a221oi_1 _5065_ (.A1(_0840_),
    .A2(_3452_),
    .B1(_3372_),
    .B2(_3456_),
    .C1(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__and4_1 _5066_ (.A(_1393_),
    .B(_1396_),
    .C(_1399_),
    .D(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__nand2_1 _5067_ (.A(_3475_),
    .B(_0708_),
    .Y(_1405_));
 sky130_fd_sc_hd__nand2_1 _5068_ (.A(_3480_),
    .B(_0334_),
    .Y(_1406_));
 sky130_fd_sc_hd__or2_1 _5069_ (.A(_3503_),
    .B(_3485_),
    .X(_1407_));
 sky130_fd_sc_hd__o2111a_1 _5070_ (.A1(_1141_),
    .A2(_3472_),
    .B1(_1405_),
    .C1(_1406_),
    .D1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__nand2_1 _5071_ (.A(_3496_),
    .B(_0329_),
    .Y(_1409_));
 sky130_fd_sc_hd__o221a_1 _5072_ (.A1(_0697_),
    .A2(_3490_),
    .B1(_3483_),
    .B2(_3493_),
    .C1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__o22ai_1 _5073_ (.A1(_3288_),
    .A2(_3502_),
    .B1(_0649_),
    .B2(_3505_),
    .Y(_1411_));
 sky130_fd_sc_hd__a22o_1 _5074_ (.A1(_3508_),
    .A2(_3246_),
    .B1(_3511_),
    .B2(_3238_),
    .X(_1412_));
 sky130_fd_sc_hd__nor2_1 _5075_ (.A(_1411_),
    .B(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__nand2_1 _5076_ (.A(_0323_),
    .B(_3287_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _5077_ (.A(_0328_),
    .B(_3512_),
    .Y(_1415_));
 sky130_fd_sc_hd__nand2_1 _5078_ (.A(_0333_),
    .B(_3275_),
    .Y(_1416_));
 sky130_fd_sc_hd__nand2_1 _5079_ (.A(_0338_),
    .B(_3509_),
    .Y(_1417_));
 sky130_fd_sc_hd__and4_1 _5080_ (.A(_1414_),
    .B(_1415_),
    .C(_1416_),
    .D(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__and4_1 _5081_ (.A(_1408_),
    .B(_1410_),
    .C(_1413_),
    .D(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__and4_1 _5082_ (.A(_1374_),
    .B(_1390_),
    .C(_1404_),
    .D(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__nor2_1 _5083_ (.A(_0394_),
    .B(_0351_),
    .Y(_1421_));
 sky130_fd_sc_hd__a22o_1 _5084_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .B1(_0356_),
    .B2(_3202_),
    .X(_1422_));
 sky130_fd_sc_hd__a211oi_1 _5085_ (.A1(_3192_),
    .A2(_0348_),
    .B1(_1421_),
    .C1(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_0370_),
    .B(_3183_),
    .Y(_1424_));
 sky130_fd_sc_hd__o21ai_1 _5087_ (.A1(_0716_),
    .A2(_0367_),
    .B1(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__a221oi_1 _5088_ (.A1(_3186_),
    .A2(_0361_),
    .B1(_3189_),
    .B2(_0364_),
    .C1(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hd__o22ai_1 _5089_ (.A1(_3488_),
    .A2(_0382_),
    .B1(_0700_),
    .B2(_0385_),
    .Y(_1427_));
 sky130_fd_sc_hd__a221oi_1 _5090_ (.A1(_0701_),
    .A2(_0376_),
    .B1(_0695_),
    .B2(_0379_),
    .C1(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__nand2_1 _5091_ (.A(_0399_),
    .B(_0634_),
    .Y(_1429_));
 sky130_fd_sc_hd__o21ai_1 _5092_ (.A1(_3491_),
    .A2(_0396_),
    .B1(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__a221oi_1 _5093_ (.A1(_3205_),
    .A2(_0390_),
    .B1(_3208_),
    .B2(_0393_),
    .C1(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__and4_1 _5094_ (.A(_1423_),
    .B(_1426_),
    .C(_1428_),
    .D(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__nand2_1 _5095_ (.A(_0412_),
    .B(_3168_),
    .Y(_1433_));
 sky130_fd_sc_hd__nand2_1 _5096_ (.A(_0417_),
    .B(_3174_),
    .Y(_1434_));
 sky130_fd_sc_hd__or2_1 _5097_ (.A(_1022_),
    .B(_0422_),
    .X(_1435_));
 sky130_fd_sc_hd__o2111a_1 _5098_ (.A1(_0349_),
    .A2(_0409_),
    .B1(_1433_),
    .C1(_1434_),
    .D1(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_0430_),
    .B(_0461_),
    .Y(_1437_));
 sky130_fd_sc_hd__nand2_1 _5100_ (.A(_0434_),
    .B(_0413_),
    .Y(_1438_));
 sky130_fd_sc_hd__or2_1 _5101_ (.A(_1175_),
    .B(_0439_),
    .X(_1439_));
 sky130_fd_sc_hd__o2111a_1 _5102_ (.A1(_0420_),
    .A2(_0427_),
    .B1(_1437_),
    .C1(_1438_),
    .D1(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__nand2_1 _5103_ (.A(_0451_),
    .B(_1039_),
    .Y(_1441_));
 sky130_fd_sc_hd__nand2_1 _5104_ (.A(_0456_),
    .B(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .Y(_1442_));
 sky130_fd_sc_hd__nand2_1 _5105_ (.A(_1441_),
    .B(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__a221oi_1 _5106_ (.A1(_0435_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0741_),
    .C1(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__nand2_1 _5107_ (.A(_0471_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _5108_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_1446_));
 sky130_fd_sc_hd__nand2_1 _5109_ (.A(_1445_),
    .B(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__a221oi_1 _5110_ (.A1(_3152_),
    .A2(_0464_),
    .B1(_3163_),
    .B2(_0468_),
    .C1(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__and4_1 _5111_ (.A(_1436_),
    .B(_1440_),
    .C(_1444_),
    .D(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(_1432_),
    .B(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _5113_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_1451_));
 sky130_fd_sc_hd__o21ai_1 _5114_ (.A1(_0920_),
    .A2(_0486_),
    .B1(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_1453_));
 sky130_fd_sc_hd__nand2_1 _5116_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_1454_));
 sky130_fd_sc_hd__nand2_1 _5117_ (.A(_1453_),
    .B(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__a221oi_1 _5118_ (.A1(_0510_),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0515_),
    .C1(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__nand2_1 _5119_ (.A(_0509_),
    .B(_0768_),
    .Y(_1457_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_0514_),
    .B(_0919_),
    .Y(_1458_));
 sky130_fd_sc_hd__and4b_1 _5121_ (.A_N(_1452_),
    .B(_1456_),
    .C(_1457_),
    .D(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__o22ai_1 _5122_ (.A1(_0772_),
    .A2(_0528_),
    .B1(_0923_),
    .B2(_0531_),
    .Y(_1460_));
 sky130_fd_sc_hd__a221oi_1 _5123_ (.A1(_0442_),
    .A2(_0521_),
    .B1(_0448_),
    .B2(_0525_),
    .C1(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__inv_2 _5124_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .Y(_1462_));
 sky130_fd_sc_hd__o22ai_1 _5125_ (.A1(_1334_),
    .A2(_0544_),
    .B1(_1462_),
    .B2(_0547_),
    .Y(_1463_));
 sky130_fd_sc_hd__a221oi_1 _5126_ (.A1(_0746_),
    .A2(_0537_),
    .B1(_0739_),
    .B2(_0541_),
    .C1(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__and3_1 _5127_ (.A(_1459_),
    .B(_1461_),
    .C(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__nand2_1 _5128_ (.A(_0563_),
    .B(_0615_),
    .Y(_1466_));
 sky130_fd_sc_hd__nand2_1 _5129_ (.A(_0568_),
    .B(_0611_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _5130_ (.A(_1466_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__a221oi_1 _5131_ (.A1(_0589_),
    .A2(_0556_),
    .B1(_0584_),
    .B2(_0560_),
    .C1(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__nand2_1 _5132_ (.A(_0583_),
    .B(_1210_),
    .Y(_1470_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(_0588_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1471_));
 sky130_fd_sc_hd__nand2_1 _5134_ (.A(_1470_),
    .B(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__a221oi_1 _5135_ (.A1(_1055_),
    .A2(_0576_),
    .B1(_1192_),
    .B2(_0580_),
    .C1(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__inv_2 _5136_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _5137_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_1475_));
 sky130_fd_sc_hd__o21ai_1 _5138_ (.A1(_1474_),
    .A2(_0603_),
    .B1(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__a221oi_1 _5139_ (.A1(_0776_),
    .A2(_0596_),
    .B1(_0927_),
    .B2(_0600_),
    .C1(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__inv_2 _5140_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_1478_));
 sky130_fd_sc_hd__o22ai_1 _5141_ (.A1(_1350_),
    .A2(_0621_),
    .B1(_1478_),
    .B2(_0624_),
    .Y(_1479_));
 sky130_fd_sc_hd__a221oi_1 _5142_ (.A1(_0781_),
    .A2(_0614_),
    .B1(_0932_),
    .B2(_0618_),
    .C1(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__and4_1 _5143_ (.A(_1469_),
    .B(_1473_),
    .C(_1477_),
    .D(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__nand2_1 _5144_ (.A(_1465_),
    .B(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__nor2_1 _5145_ (.A(_1450_),
    .B(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__nand2_1 _5146_ (.A(_0633_),
    .B(_3476_),
    .Y(_1484_));
 sky130_fd_sc_hd__nand3_2 _5147_ (.A(_1420_),
    .B(_1483_),
    .C(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__nor2_1 _5148_ (.A(_3212_),
    .B(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__nor2_1 _5149_ (.A(_1359_),
    .B(_1486_),
    .Y(_0291_));
 sky130_fd_sc_hd__o21ai_1 _5150_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B1(_3161_),
    .Y(_1487_));
 sky130_fd_sc_hd__nand2_1 _5151_ (.A(_3237_),
    .B(_3271_),
    .Y(_1488_));
 sky130_fd_sc_hd__nand2_1 _5152_ (.A(_3245_),
    .B(_3306_),
    .Y(_1489_));
 sky130_fd_sc_hd__nand2_1 _5153_ (.A(_1488_),
    .B(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__a221oi_1 _5154_ (.A1(_3264_),
    .A2(_3223_),
    .B1(_3250_),
    .B2(_3229_),
    .C1(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_3263_),
    .B(_0991_),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_1 _5156_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .Y(_1493_));
 sky130_fd_sc_hd__nand2_1 _5157_ (.A(_1492_),
    .B(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__a221oi_1 _5158_ (.A1(_1130_),
    .A2(_3254_),
    .B1(_3395_),
    .B2(_3258_),
    .C1(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_3295_),
    .B(_3300_),
    .Y(_1496_));
 sky130_fd_sc_hd__o21ai_1 _5160_ (.A1(_3315_),
    .A2(_3291_),
    .B1(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__a221oi_1 _5161_ (.A1(_3224_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_0639_),
    .C1(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__inv_2 _5162_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_1499_));
 sky130_fd_sc_hd__o22ai_1 _5163_ (.A1(_1371_),
    .A2(_3314_),
    .B1(_1499_),
    .B2(_3318_),
    .Y(_1500_));
 sky130_fd_sc_hd__a221oi_1 _5164_ (.A1(_3439_),
    .A2(_3305_),
    .B1(_0683_),
    .B2(_3310_),
    .C1(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__and4_1 _5165_ (.A(_1491_),
    .B(_1495_),
    .C(_1498_),
    .D(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__nand2_1 _5166_ (.A(_3335_),
    .B(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_1503_));
 sky130_fd_sc_hd__o21ai_1 _5167_ (.A1(_1474_),
    .A2(_3332_),
    .B1(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__a221oi_1 _5168_ (.A1(_0597_),
    .A2(_3326_),
    .B1(_0569_),
    .B2(_3330_),
    .C1(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__inv_2 _5169_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_1506_));
 sky130_fd_sc_hd__nand2_1 _5170_ (.A(_3353_),
    .B(_3327_),
    .Y(_1507_));
 sky130_fd_sc_hd__o21ai_1 _5171_ (.A1(_1506_),
    .A2(_3350_),
    .B1(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__a221oi_1 _5172_ (.A1(_3380_),
    .A2(_3343_),
    .B1(_3322_),
    .B2(_3347_),
    .C1(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(_3371_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1510_));
 sky130_fd_sc_hd__o21ai_1 _5174_ (.A1(_3348_),
    .A2(_3368_),
    .B1(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__a221oi_1 _5175_ (.A1(_0972_),
    .A2(_3361_),
    .B1(_3376_),
    .B2(_3365_),
    .C1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand2_1 _5176_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_1513_));
 sky130_fd_sc_hd__nand2_1 _5177_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_1514_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(_1513_),
    .B(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__a221oi_1 _5179_ (.A1(_0607_),
    .A2(_3379_),
    .B1(_0593_),
    .B2(_3383_),
    .C1(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__and4_1 _5180_ (.A(_1505_),
    .B(_1509_),
    .C(_1512_),
    .D(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__inv_2 _5181_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1518_));
 sky130_fd_sc_hd__o22ai_1 _5182_ (.A1(_1391_),
    .A2(_3408_),
    .B1(_1518_),
    .B2(_3411_),
    .Y(_1519_));
 sky130_fd_sc_hd__a221oi_1 _5183_ (.A1(_3418_),
    .A2(_3401_),
    .B1(_3428_),
    .B2(_3405_),
    .C1(_1519_),
    .Y(_1520_));
 sky130_fd_sc_hd__nand2_1 _5184_ (.A(_3427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1521_));
 sky130_fd_sc_hd__o21ai_1 _5185_ (.A1(_1382_),
    .A2(_3424_),
    .B1(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__a221oi_1 _5186_ (.A1(_3362_),
    .A2(_3417_),
    .B1(_3340_),
    .B2(_3421_),
    .C1(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__nand2_1 _5187_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .Y(_1524_));
 sky130_fd_sc_hd__o21ai_1 _5188_ (.A1(_1124_),
    .A2(_3442_),
    .B1(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__a221oi_1 _5189_ (.A1(_3402_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_0675_),
    .C1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _5190_ (.A(_3459_),
    .B(_0840_),
    .Y(_1527_));
 sky130_fd_sc_hd__nand2_1 _5191_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .Y(_1528_));
 sky130_fd_sc_hd__nand2_1 _5192_ (.A(_1527_),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__a221oi_1 _5193_ (.A1(_3372_),
    .A2(_3452_),
    .B1(_3358_),
    .B2(_3456_),
    .C1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__and4_1 _5194_ (.A(_1520_),
    .B(_1523_),
    .C(_1526_),
    .D(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__nand2_1 _5195_ (.A(_3475_),
    .B(_0865_),
    .Y(_1532_));
 sky130_fd_sc_hd__nand2_1 _5196_ (.A(_3480_),
    .B(_0324_),
    .Y(_1533_));
 sky130_fd_sc_hd__or2_1 _5197_ (.A(_0704_),
    .B(_3485_),
    .X(_1534_));
 sky130_fd_sc_hd__o2111a_1 _5198_ (.A1(_3500_),
    .A2(_3472_),
    .B1(_1532_),
    .C1(_1533_),
    .D1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__nand2_1 _5199_ (.A(_3496_),
    .B(_0334_),
    .Y(_1536_));
 sky130_fd_sc_hd__o221a_1 _5200_ (.A1(_0855_),
    .A2(_3490_),
    .B1(_0697_),
    .B2(_3493_),
    .C1(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__o22ai_1 _5201_ (.A1(_0649_),
    .A2(_3502_),
    .B1(_0810_),
    .B2(_3505_),
    .Y(_1538_));
 sky130_fd_sc_hd__a22o_1 _5202_ (.A1(_3508_),
    .A2(_3238_),
    .B1(_3511_),
    .B2(_3213_),
    .X(_1539_));
 sky130_fd_sc_hd__nor2_1 _5203_ (.A(_1538_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__nand2_1 _5204_ (.A(_0323_),
    .B(_0648_),
    .Y(_1541_));
 sky130_fd_sc_hd__nand2_1 _5205_ (.A(_0328_),
    .B(_3275_),
    .Y(_1542_));
 sky130_fd_sc_hd__nand2_1 _5206_ (.A(_0333_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _5207_ (.A(_0338_),
    .B(_3512_),
    .Y(_1544_));
 sky130_fd_sc_hd__and4_1 _5208_ (.A(_1541_),
    .B(_1542_),
    .C(_1543_),
    .D(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__and4_1 _5209_ (.A(_1535_),
    .B(_1537_),
    .C(_1540_),
    .D(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__and4_1 _5210_ (.A(_1502_),
    .B(_1517_),
    .C(_1531_),
    .D(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__nor2_1 _5211_ (.A(_0380_),
    .B(_0351_),
    .Y(_1548_));
 sky130_fd_sc_hd__a22o_1 _5212_ (.A1(_0354_),
    .A2(_3202_),
    .B1(_0356_),
    .B2(_3205_),
    .X(_1549_));
 sky130_fd_sc_hd__a211oi_1 _5213_ (.A1(_3195_),
    .A2(_0348_),
    .B1(_1548_),
    .C1(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__nand2_1 _5214_ (.A(_0370_),
    .B(_3186_),
    .Y(_1551_));
 sky130_fd_sc_hd__o21ai_1 _5215_ (.A1(_0873_),
    .A2(_0367_),
    .B1(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__a221oi_1 _5216_ (.A1(_3189_),
    .A2(_0361_),
    .B1(_3192_),
    .B2(_0364_),
    .C1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__o22ai_1 _5217_ (.A1(_0700_),
    .A2(_0382_),
    .B1(_0858_),
    .B2(_0385_),
    .Y(_1554_));
 sky130_fd_sc_hd__a221oi_1 _5218_ (.A1(_0695_),
    .A2(_0376_),
    .B1(_3476_),
    .B2(_0379_),
    .C1(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_1 _5219_ (.A(_0399_),
    .B(_0796_),
    .Y(_1556_));
 sky130_fd_sc_hd__o21ai_1 _5220_ (.A1(_3488_),
    .A2(_0396_),
    .B1(_1556_),
    .Y(_1557_));
 sky130_fd_sc_hd__a221oi_1 _5221_ (.A1(_3208_),
    .A2(_0390_),
    .B1(_0634_),
    .B2(_0393_),
    .C1(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__and4_1 _5222_ (.A(_1550_),
    .B(_1553_),
    .C(_1555_),
    .D(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__nand2_1 _5223_ (.A(_0412_),
    .B(_3171_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2_1 _5224_ (.A(_0417_),
    .B(_3177_),
    .Y(_1561_));
 sky130_fd_sc_hd__or2_1 _5225_ (.A(_1161_),
    .B(_0422_),
    .X(_1562_));
 sky130_fd_sc_hd__o2111a_1 _5226_ (.A1(_0716_),
    .A2(_0409_),
    .B1(_1560_),
    .C1(_1561_),
    .D1(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__nand2_1 _5227_ (.A(_0430_),
    .B(_0465_),
    .Y(_1564_));
 sky130_fd_sc_hd__nand2_1 _5228_ (.A(_0434_),
    .B(_0731_),
    .Y(_1565_));
 sky130_fd_sc_hd__or2_1 _5229_ (.A(_1308_),
    .B(_0439_),
    .X(_1566_));
 sky130_fd_sc_hd__o2111a_1 _5230_ (.A1(_0735_),
    .A2(_0427_),
    .B1(_1564_),
    .C1(_1565_),
    .D1(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__nand2_1 _5231_ (.A(_0451_),
    .B(_0461_),
    .Y(_1568_));
 sky130_fd_sc_hd__nand2_1 _5232_ (.A(_0456_),
    .B(_1039_),
    .Y(_1569_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_1568_),
    .B(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__a221oi_1 _5234_ (.A1(_0741_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0894_),
    .C1(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_1 _5235_ (.A(_0471_),
    .B(_3152_),
    .Y(_1572_));
 sky130_fd_sc_hd__nand2_1 _5236_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2_1 _5237_ (.A(_1572_),
    .B(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__a221oi_1 _5238_ (.A1(_3163_),
    .A2(_0464_),
    .B1(_3168_),
    .B2(_0468_),
    .C1(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hd__and4_1 _5239_ (.A(_1563_),
    .B(_1567_),
    .C(_1571_),
    .D(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__nand2_1 _5240_ (.A(_1559_),
    .B(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__nand2_1 _5241_ (.A(_0489_),
    .B(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_1578_));
 sky130_fd_sc_hd__o21ai_1 _5242_ (.A1(_0542_),
    .A2(_0486_),
    .B1(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_1580_));
 sky130_fd_sc_hd__nand2_1 _5244_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_1581_));
 sky130_fd_sc_hd__nand2_1 _5245_ (.A(_1580_),
    .B(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__a221oi_1 _5246_ (.A1(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0765_),
    .C1(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(_0509_),
    .B(_0919_),
    .Y(_1584_));
 sky130_fd_sc_hd__nand2_1 _5248_ (.A(_0514_),
    .B(_0534_),
    .Y(_1585_));
 sky130_fd_sc_hd__and4b_1 _5249_ (.A_N(_1579_),
    .B(_1583_),
    .C(_1584_),
    .D(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__o22ai_1 _5250_ (.A1(_0923_),
    .A2(_0528_),
    .B1(_1065_),
    .B2(_0531_),
    .Y(_1587_));
 sky130_fd_sc_hd__a221oi_1 _5251_ (.A1(_0448_),
    .A2(_0521_),
    .B1(_0457_),
    .B2(_0525_),
    .C1(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__inv_2 _5252_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_1589_));
 sky130_fd_sc_hd__o22ai_1 _5253_ (.A1(_1462_),
    .A2(_0544_),
    .B1(_1589_),
    .B2(_0547_),
    .Y(_1590_));
 sky130_fd_sc_hd__a221oi_1 _5254_ (.A1(_0739_),
    .A2(_0537_),
    .B1(_0435_),
    .B2(_0541_),
    .C1(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__and3_1 _5255_ (.A(_1586_),
    .B(_1588_),
    .C(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(_0563_),
    .B(_0589_),
    .Y(_1593_));
 sky130_fd_sc_hd__nand2_1 _5257_ (.A(_0568_),
    .B(_0615_),
    .Y(_1594_));
 sky130_fd_sc_hd__nand2_1 _5258_ (.A(_1593_),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__a221oi_1 _5259_ (.A1(_0584_),
    .A2(_0556_),
    .B1(_0573_),
    .B2(_0560_),
    .C1(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _5260_ (.A(_0583_),
    .B(_1055_),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _5261_ (.A(_0588_),
    .B(_1210_),
    .Y(_1598_));
 sky130_fd_sc_hd__nand2_1 _5262_ (.A(_1597_),
    .B(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__a221oi_1 _5263_ (.A1(_1192_),
    .A2(_0576_),
    .B1(_0510_),
    .B2(_0580_),
    .C1(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__inv_2 _5264_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_1601_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_1602_));
 sky130_fd_sc_hd__o21ai_1 _5266_ (.A1(_1601_),
    .A2(_0603_),
    .B1(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__a221oi_1 _5267_ (.A1(_0927_),
    .A2(_0596_),
    .B1(_0611_),
    .B2(_0600_),
    .C1(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__inv_2 _5268_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_1605_));
 sky130_fd_sc_hd__o22ai_1 _5269_ (.A1(_1478_),
    .A2(_0621_),
    .B1(_1605_),
    .B2(_0624_),
    .Y(_1606_));
 sky130_fd_sc_hd__a221oi_1 _5270_ (.A1(_0932_),
    .A2(_0614_),
    .B1(_1073_),
    .B2(_0618_),
    .C1(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__and4_1 _5271_ (.A(_1596_),
    .B(_1600_),
    .C(_1604_),
    .D(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__nand2_1 _5272_ (.A(_1592_),
    .B(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__nor2_1 _5273_ (.A(_1577_),
    .B(_1609_),
    .Y(_1610_));
 sky130_fd_sc_hd__nand2_1 _5274_ (.A(_0633_),
    .B(_3482_),
    .Y(_1611_));
 sky130_fd_sc_hd__nand3_2 _5275_ (.A(_1547_),
    .B(_1610_),
    .C(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__nor2_1 _5276_ (.A(_3212_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__nor2_1 _5277_ (.A(_1487_),
    .B(_1613_),
    .Y(_0290_));
 sky130_fd_sc_hd__o21ai_1 _5278_ (.A1(_3151_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B1(_3161_),
    .Y(_1614_));
 sky130_fd_sc_hd__nand2_1 _5279_ (.A(_3237_),
    .B(_3264_),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2_1 _5280_ (.A(_3245_),
    .B(_3271_),
    .Y(_1616_));
 sky130_fd_sc_hd__nand2_1 _5281_ (.A(_1615_),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__a221oi_1 _5282_ (.A1(_3250_),
    .A2(_3223_),
    .B1(_3255_),
    .B2(_3229_),
    .C1(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__nand2_1 _5283_ (.A(_3263_),
    .B(_1130_),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2_1 _5284_ (.A(_3270_),
    .B(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .Y(_1620_));
 sky130_fd_sc_hd__nand2_1 _5285_ (.A(_1619_),
    .B(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__a221oi_1 _5286_ (.A1(_3395_),
    .A2(_3254_),
    .B1(_3402_),
    .B2(_3258_),
    .C1(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__nand2_1 _5287_ (.A(_3295_),
    .B(_3306_),
    .Y(_1623_));
 sky130_fd_sc_hd__o21ai_1 _5288_ (.A1(_0653_),
    .A2(_3291_),
    .B1(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__a221oi_1 _5289_ (.A1(_0639_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_0801_),
    .C1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__inv_2 _5290_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_1626_));
 sky130_fd_sc_hd__o22ai_1 _5291_ (.A1(_1499_),
    .A2(_3314_),
    .B1(_1626_),
    .B2(_3318_),
    .Y(_1627_));
 sky130_fd_sc_hd__a221oi_1 _5292_ (.A1(_0683_),
    .A2(_3305_),
    .B1(_0844_),
    .B2(_3310_),
    .C1(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__and4_1 _5293_ (.A(_1618_),
    .B(_1622_),
    .C(_1625_),
    .D(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__nand2_1 _5294_ (.A(_3335_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1630_));
 sky130_fd_sc_hd__o21ai_1 _5295_ (.A1(_1601_),
    .A2(_3332_),
    .B1(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__a221oi_1 _5296_ (.A1(_0569_),
    .A2(_3326_),
    .B1(_0564_),
    .B2(_3330_),
    .C1(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__nand2_1 _5297_ (.A(_3353_),
    .B(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_1633_));
 sky130_fd_sc_hd__o21ai_1 _5298_ (.A1(_3331_),
    .A2(_3350_),
    .B1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__a221oi_1 _5299_ (.A1(_3322_),
    .A2(_3343_),
    .B1(_3327_),
    .B2(_3347_),
    .C1(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(_3371_),
    .B(_0972_),
    .Y(_1636_));
 sky130_fd_sc_hd__o21ai_1 _5301_ (.A1(_0661_),
    .A2(_3368_),
    .B1(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__a221oi_1 _5302_ (.A1(_3376_),
    .A2(_3361_),
    .B1(_3380_),
    .B2(_3365_),
    .C1(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__nand2_1 _5303_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_1639_));
 sky130_fd_sc_hd__nand2_1 _5304_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_1640_));
 sky130_fd_sc_hd__nand2_1 _5305_ (.A(_1639_),
    .B(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__a221oi_1 _5306_ (.A1(_0593_),
    .A2(_3379_),
    .B1(_0597_),
    .B2(_3383_),
    .C1(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__and4_1 _5307_ (.A(_1632_),
    .B(_1635_),
    .C(_1638_),
    .D(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__inv_2 _5308_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1644_));
 sky130_fd_sc_hd__o22ai_1 _5309_ (.A1(_1518_),
    .A2(_3408_),
    .B1(_1644_),
    .B2(_3411_),
    .Y(_1645_));
 sky130_fd_sc_hd__a221oi_1 _5310_ (.A1(_3428_),
    .A2(_3401_),
    .B1(_0679_),
    .B2(_3405_),
    .C1(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__nand2_1 _5311_ (.A(_3427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1647_));
 sky130_fd_sc_hd__o21ai_1 _5312_ (.A1(_3348_),
    .A2(_3424_),
    .B1(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__a221oi_1 _5313_ (.A1(_3340_),
    .A2(_3417_),
    .B1(_3344_),
    .B2(_3421_),
    .C1(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__nand2_1 _5314_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .Y(_1650_));
 sky130_fd_sc_hd__o21ai_1 _5315_ (.A1(_1261_),
    .A2(_3442_),
    .B1(_1650_),
    .Y(_1651_));
 sky130_fd_sc_hd__a221oi_1 _5316_ (.A1(_0675_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_0836_),
    .C1(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__nand2_1 _5317_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_1653_));
 sky130_fd_sc_hd__nand2_1 _5318_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .Y(_1654_));
 sky130_fd_sc_hd__nand2_1 _5319_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__a221oi_1 _5320_ (.A1(_3358_),
    .A2(_3452_),
    .B1(_3362_),
    .B2(_3456_),
    .C1(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__and4_1 _5321_ (.A(_1646_),
    .B(_1649_),
    .C(_1652_),
    .D(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__nand2_1 _5322_ (.A(_3475_),
    .B(_3509_),
    .Y(_1658_));
 sky130_fd_sc_hd__nand2_1 _5323_ (.A(_3480_),
    .B(_0708_),
    .Y(_1659_));
 sky130_fd_sc_hd__or2_1 _5324_ (.A(_0861_),
    .B(_3485_),
    .X(_1660_));
 sky130_fd_sc_hd__o2111a_1 _5325_ (.A1(_3503_),
    .A2(_3472_),
    .B1(_1658_),
    .C1(_1659_),
    .D1(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__nand2_1 _5326_ (.A(_3496_),
    .B(_0324_),
    .Y(_1662_));
 sky130_fd_sc_hd__o221a_1 _5327_ (.A1(_1002_),
    .A2(_3490_),
    .B1(_0855_),
    .B2(_3493_),
    .C1(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__o22ai_1 _5328_ (.A1(_0810_),
    .A2(_3502_),
    .B1(_0960_),
    .B2(_3505_),
    .Y(_1664_));
 sky130_fd_sc_hd__a22o_1 _5329_ (.A1(_3508_),
    .A2(_3213_),
    .B1(_3511_),
    .B2(_3224_),
    .X(_1665_));
 sky130_fd_sc_hd__nor2_1 _5330_ (.A(_1664_),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__nand2_1 _5331_ (.A(_0323_),
    .B(_3296_),
    .Y(_1667_));
 sky130_fd_sc_hd__nand2_1 _5332_ (.A(_0328_),
    .B(_3287_),
    .Y(_1668_));
 sky130_fd_sc_hd__nand2_1 _5333_ (.A(_0333_),
    .B(_0648_),
    .Y(_1669_));
 sky130_fd_sc_hd__nand2_1 _5334_ (.A(_0338_),
    .B(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .Y(_1670_));
 sky130_fd_sc_hd__and4_1 _5335_ (.A(_1667_),
    .B(_1668_),
    .C(_1669_),
    .D(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__and4_1 _5336_ (.A(_1661_),
    .B(_1663_),
    .C(_1666_),
    .D(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__and4_1 _5337_ (.A(_1629_),
    .B(_1643_),
    .C(_1657_),
    .D(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__nor2_1 _5338_ (.A(_0383_),
    .B(_0351_),
    .Y(_1674_));
 sky130_fd_sc_hd__a22o_1 _5339_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .B1(_0356_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_1675_));
 sky130_fd_sc_hd__a211oi_1 _5340_ (.A1(_3199_),
    .A2(_0348_),
    .B1(_1674_),
    .C1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand2_1 _5341_ (.A(_0370_),
    .B(_3189_),
    .Y(_1677_));
 sky130_fd_sc_hd__o21ai_1 _5342_ (.A1(_1018_),
    .A2(_0367_),
    .B1(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__a221oi_1 _5343_ (.A1(_3192_),
    .A2(_0361_),
    .B1(_3195_),
    .B2(_0364_),
    .C1(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__o22ai_1 _5344_ (.A1(_0858_),
    .A2(_0382_),
    .B1(_3468_),
    .B2(_0385_),
    .Y(_1680_));
 sky130_fd_sc_hd__a221oi_1 _5345_ (.A1(_3476_),
    .A2(_0376_),
    .B1(_3482_),
    .B2(_0379_),
    .C1(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__nand2_1 _5346_ (.A(_0399_),
    .B(_0947_),
    .Y(_1682_));
 sky130_fd_sc_hd__o21ai_1 _5347_ (.A1(_0700_),
    .A2(_0396_),
    .B1(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__a221oi_1 _5348_ (.A1(_0634_),
    .A2(_0390_),
    .B1(_0796_),
    .B2(_0393_),
    .C1(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__and4_1 _5349_ (.A(_1676_),
    .B(_1679_),
    .C(_1681_),
    .D(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_1 _5350_ (.A(_0412_),
    .B(_3174_),
    .Y(_1686_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(_0417_),
    .B(_3180_),
    .Y(_1687_));
 sky130_fd_sc_hd__or2_1 _5352_ (.A(_0349_),
    .B(_0422_),
    .X(_1688_));
 sky130_fd_sc_hd__o2111a_1 _5353_ (.A1(_0873_),
    .A2(_0409_),
    .B1(_1686_),
    .C1(_1687_),
    .D1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__nand2_1 _5354_ (.A(_0430_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1690_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_0434_),
    .B(_0418_),
    .Y(_1691_));
 sky130_fd_sc_hd__or2_1 _5356_ (.A(_0420_),
    .B(_0439_),
    .X(_1692_));
 sky130_fd_sc_hd__o2111a_1 _5357_ (.A1(_0404_),
    .A2(_0427_),
    .B1(_1690_),
    .C1(_1691_),
    .D1(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__nand2_1 _5358_ (.A(_0451_),
    .B(_0465_),
    .Y(_1694_));
 sky130_fd_sc_hd__nand2_1 _5359_ (.A(_0456_),
    .B(_0461_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand2_1 _5360_ (.A(_1694_),
    .B(_1695_),
    .Y(_1696_));
 sky130_fd_sc_hd__a221oi_2 _5361_ (.A1(_0894_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_1039_),
    .C1(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(_0471_),
    .B(_3163_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_1 _5363_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_1 _5364_ (.A(_1698_),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__a221oi_1 _5365_ (.A1(_3168_),
    .A2(_0464_),
    .B1(_3171_),
    .B2(_0468_),
    .C1(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__and4_1 _5366_ (.A(_1689_),
    .B(_1693_),
    .C(_1697_),
    .D(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__nand2_1 _5367_ (.A(_1685_),
    .B(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__nand2_1 _5368_ (.A(_0489_),
    .B(_0768_),
    .Y(_1704_));
 sky130_fd_sc_hd__o21ai_1 _5369_ (.A1(_0545_),
    .A2(_0486_),
    .B1(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_1706_));
 sky130_fd_sc_hd__nand2_1 _5371_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_1707_));
 sky130_fd_sc_hd__nand2_1 _5372_ (.A(_1706_),
    .B(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__a221oi_1 _5373_ (.A1(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0916_),
    .C1(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand2_1 _5374_ (.A(_0509_),
    .B(_0534_),
    .Y(_1710_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(_0514_),
    .B(_0538_),
    .Y(_1711_));
 sky130_fd_sc_hd__and4b_1 _5376_ (.A_N(_1705_),
    .B(_1709_),
    .C(_1710_),
    .D(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__o22ai_1 _5377_ (.A1(_1065_),
    .A2(_0528_),
    .B1(_1202_),
    .B2(_0531_),
    .Y(_1713_));
 sky130_fd_sc_hd__a221oi_1 _5378_ (.A1(_0457_),
    .A2(_0521_),
    .B1(_0452_),
    .B2(_0525_),
    .C1(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__o22ai_1 _5379_ (.A1(_1589_),
    .A2(_0544_),
    .B1(_0437_),
    .B2(_0547_),
    .Y(_1715_));
 sky130_fd_sc_hd__a221oi_1 _5380_ (.A1(_0435_),
    .A2(_0537_),
    .B1(_0741_),
    .B2(_0541_),
    .C1(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__and3_1 _5381_ (.A(_1712_),
    .B(_1714_),
    .C(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__nand2_1 _5382_ (.A(_0563_),
    .B(_0584_),
    .Y(_1718_));
 sky130_fd_sc_hd__nand2_1 _5383_ (.A(_0568_),
    .B(_0589_),
    .Y(_1719_));
 sky130_fd_sc_hd__nand2_1 _5384_ (.A(_1718_),
    .B(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__a221oi_1 _5385_ (.A1(_0573_),
    .A2(_0556_),
    .B1(_0577_),
    .B2(_0560_),
    .C1(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_1 _5386_ (.A(_0583_),
    .B(_1192_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand2_1 _5387_ (.A(_0588_),
    .B(_1055_),
    .Y(_1723_));
 sky130_fd_sc_hd__nand2_1 _5388_ (.A(_1722_),
    .B(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__a221oi_1 _5389_ (.A1(_0510_),
    .A2(_0576_),
    .B1(_0515_),
    .B2(_0580_),
    .C1(_1724_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_1726_));
 sky130_fd_sc_hd__o21ai_1 _5391_ (.A1(_0619_),
    .A2(_0603_),
    .B1(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__a221oi_1 _5392_ (.A1(_0611_),
    .A2(_0596_),
    .B1(_0615_),
    .B2(_0600_),
    .C1(_1727_),
    .Y(_1728_));
 sky130_fd_sc_hd__inv_2 _5393_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1729_));
 sky130_fd_sc_hd__o22ai_1 _5394_ (.A1(_1605_),
    .A2(_0621_),
    .B1(_1729_),
    .B2(_0624_),
    .Y(_1730_));
 sky130_fd_sc_hd__a221oi_1 _5395_ (.A1(_1073_),
    .A2(_0614_),
    .B1(_1210_),
    .B2(_0618_),
    .C1(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__and4_1 _5396_ (.A(_1721_),
    .B(_1725_),
    .C(_1728_),
    .D(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__nand2_1 _5397_ (.A(_1717_),
    .B(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__nor2_1 _5398_ (.A(_1703_),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _5399_ (.A(_0633_),
    .B(_0339_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand3_1 _5400_ (.A(_1673_),
    .B(_1734_),
    .C(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__nor2_1 _5401_ (.A(_3212_),
    .B(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__nor2_1 _5402_ (.A(_1614_),
    .B(_1737_),
    .Y(_0289_));
 sky130_fd_sc_hd__o21ai_1 _5403_ (.A1(_3150_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B1(_3161_),
    .Y(_1738_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(_3237_),
    .B(_3250_),
    .Y(_1739_));
 sky130_fd_sc_hd__nand2_1 _5405_ (.A(_3245_),
    .B(_3264_),
    .Y(_1740_));
 sky130_fd_sc_hd__nand2_1 _5406_ (.A(_1739_),
    .B(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hd__a221oi_2 _5407_ (.A1(_3255_),
    .A2(_3223_),
    .B1(_3432_),
    .B2(_3229_),
    .C1(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_3263_),
    .B(_3395_),
    .Y(_1743_));
 sky130_fd_sc_hd__nand2_1 _5409_ (.A(_3270_),
    .B(_1130_),
    .Y(_1744_));
 sky130_fd_sc_hd__nand2_1 _5410_ (.A(_1743_),
    .B(_1744_),
    .Y(_1745_));
 sky130_fd_sc_hd__a221oi_1 _5411_ (.A1(_3402_),
    .A2(_3254_),
    .B1(_0675_),
    .B2(_3258_),
    .C1(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5412_ (.A(_3295_),
    .B(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .Y(_1747_));
 sky130_fd_sc_hd__o21ai_1 _5413_ (.A1(_0814_),
    .A2(_3291_),
    .B1(_1747_),
    .Y(_1748_));
 sky130_fd_sc_hd__a221oi_1 _5414_ (.A1(_0801_),
    .A2(_3281_),
    .B1(_3286_),
    .B2(_3300_),
    .C1(_1748_),
    .Y(_1749_));
 sky130_fd_sc_hd__o22ai_1 _5415_ (.A1(_1626_),
    .A2(_3314_),
    .B1(_3440_),
    .B2(_3318_),
    .Y(_1750_));
 sky130_fd_sc_hd__a221oi_1 _5416_ (.A1(_0844_),
    .A2(_3305_),
    .B1(_0991_),
    .B2(_3310_),
    .C1(_1750_),
    .Y(_1751_));
 sky130_fd_sc_hd__and4_1 _5417_ (.A(_1742_),
    .B(_1746_),
    .C(_1749_),
    .D(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__nand2_1 _5418_ (.A(_3335_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_1753_));
 sky130_fd_sc_hd__o21ai_1 _5419_ (.A1(_0619_),
    .A2(_3332_),
    .B1(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__a221oi_1 _5420_ (.A1(_0564_),
    .A2(_3326_),
    .B1(_0551_),
    .B2(_3330_),
    .C1(_1754_),
    .Y(_1755_));
 sky130_fd_sc_hd__nand2_1 _5421_ (.A(_3353_),
    .B(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_1756_));
 sky130_fd_sc_hd__o21ai_1 _5422_ (.A1(_0601_),
    .A2(_3350_),
    .B1(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__a221oi_1 _5423_ (.A1(_3327_),
    .A2(_3343_),
    .B1(_3336_),
    .B2(_3347_),
    .C1(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__nand2_1 _5424_ (.A(_3371_),
    .B(_3376_),
    .Y(_1759_));
 sky130_fd_sc_hd__o21ai_1 _5425_ (.A1(_0822_),
    .A2(_3368_),
    .B1(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hd__a221oi_1 _5426_ (.A1(_3380_),
    .A2(_3361_),
    .B1(_3322_),
    .B2(_3365_),
    .C1(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_3386_),
    .B(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_1762_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_3390_),
    .B(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_1763_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1762_),
    .B(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__a221oi_2 _5430_ (.A1(_0597_),
    .A2(_3379_),
    .B1(_0569_),
    .B2(_3383_),
    .C1(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__and4_1 _5431_ (.A(_1755_),
    .B(_1758_),
    .C(_1761_),
    .D(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__inv_2 _5432_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1767_));
 sky130_fd_sc_hd__o22ai_1 _5433_ (.A1(_1644_),
    .A2(_3408_),
    .B1(_1767_),
    .B2(_3411_),
    .Y(_1768_));
 sky130_fd_sc_hd__a221oi_1 _5434_ (.A1(_0679_),
    .A2(_3401_),
    .B1(_0840_),
    .B2(_3405_),
    .C1(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__nand2_1 _5435_ (.A(_3427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1770_));
 sky130_fd_sc_hd__o21ai_1 _5436_ (.A1(_0661_),
    .A2(_3424_),
    .B1(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__a221oi_1 _5437_ (.A1(_3344_),
    .A2(_3417_),
    .B1(_3354_),
    .B2(_3421_),
    .C1(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(_3445_),
    .B(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .Y(_1773_));
 sky130_fd_sc_hd__o21ai_1 _5439_ (.A1(_1391_),
    .A2(_3442_),
    .B1(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__a221oi_1 _5440_ (.A1(_0836_),
    .A2(_3435_),
    .B1(_3438_),
    .B2(_3449_),
    .C1(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(_3459_),
    .B(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_1776_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_3463_),
    .B(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .Y(_1777_));
 sky130_fd_sc_hd__nand2_1 _5443_ (.A(_1776_),
    .B(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__a221oi_1 _5444_ (.A1(_3362_),
    .A2(_3452_),
    .B1(_3340_),
    .B2(_3456_),
    .C1(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__and4_1 _5445_ (.A(_1769_),
    .B(_1772_),
    .C(_1775_),
    .D(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__nand2_1 _5446_ (.A(_3475_),
    .B(_3512_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_1 _5447_ (.A(_3480_),
    .B(_0865_),
    .Y(_1782_));
 sky130_fd_sc_hd__or2_1 _5448_ (.A(_1007_),
    .B(_3485_),
    .X(_1783_));
 sky130_fd_sc_hd__o2111a_1 _5449_ (.A1(_0704_),
    .A2(_3472_),
    .B1(_1781_),
    .C1(_1782_),
    .D1(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__nand2_1 _5450_ (.A(_3496_),
    .B(_0708_),
    .Y(_1785_));
 sky130_fd_sc_hd__o221a_1 _5451_ (.A1(_1141_),
    .A2(_3490_),
    .B1(_1002_),
    .B2(_3493_),
    .C1(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__o22ai_1 _5452_ (.A1(_0960_),
    .A2(_3502_),
    .B1(_1100_),
    .B2(_3505_),
    .Y(_1787_));
 sky130_fd_sc_hd__a22o_1 _5453_ (.A1(_3508_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .B1(_3511_),
    .B2(_0639_),
    .X(_1788_));
 sky130_fd_sc_hd__nor2_1 _5454_ (.A(_1787_),
    .B(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__nand2_1 _5455_ (.A(_0323_),
    .B(_3246_),
    .Y(_1790_));
 sky130_fd_sc_hd__nand2_1 _5456_ (.A(_0328_),
    .B(_0648_),
    .Y(_1791_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(_0333_),
    .B(_3296_),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_0338_),
    .B(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .Y(_1793_));
 sky130_fd_sc_hd__and4_1 _5459_ (.A(_1790_),
    .B(_1791_),
    .C(_1792_),
    .D(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__and4_1 _5460_ (.A(_1784_),
    .B(_1786_),
    .C(_1789_),
    .D(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__and4_1 _5461_ (.A(_1752_),
    .B(_1766_),
    .C(_1780_),
    .D(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__nor2_1 _5462_ (.A(_0724_),
    .B(_0351_),
    .Y(_1797_));
 sky130_fd_sc_hd__a22o_1 _5463_ (.A1(_0354_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .B1(_0356_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_1798_));
 sky130_fd_sc_hd__a211oi_1 _5464_ (.A1(_3202_),
    .A2(_0348_),
    .B1(_1797_),
    .C1(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_0370_),
    .B(_3192_),
    .Y(_1800_));
 sky130_fd_sc_hd__o21ai_1 _5466_ (.A1(_1157_),
    .A2(_0367_),
    .B1(_1800_),
    .Y(_1801_));
 sky130_fd_sc_hd__a221oi_1 _5467_ (.A1(_3195_),
    .A2(_0361_),
    .B1(_3199_),
    .B2(_0364_),
    .C1(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__o22ai_1 _5468_ (.A1(_3468_),
    .A2(_0382_),
    .B1(_0693_),
    .B2(_0385_),
    .Y(_1803_));
 sky130_fd_sc_hd__a221oi_1 _5469_ (.A1(_3482_),
    .A2(_0376_),
    .B1(_0339_),
    .B2(_0379_),
    .C1(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__nand2_1 _5470_ (.A(_0399_),
    .B(_3497_),
    .Y(_1805_));
 sky130_fd_sc_hd__o21ai_1 _5471_ (.A1(_0858_),
    .A2(_0396_),
    .B1(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__a221oi_1 _5472_ (.A1(_0796_),
    .A2(_0390_),
    .B1(_0947_),
    .B2(_0393_),
    .C1(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__and4_1 _5473_ (.A(_1799_),
    .B(_1802_),
    .C(_1804_),
    .D(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__nand2_1 _5474_ (.A(_0412_),
    .B(_3177_),
    .Y(_1809_));
 sky130_fd_sc_hd__nand2_1 _5475_ (.A(_0417_),
    .B(_3183_),
    .Y(_1810_));
 sky130_fd_sc_hd__or2_1 _5476_ (.A(_0716_),
    .B(_0422_),
    .X(_1811_));
 sky130_fd_sc_hd__o2111a_1 _5477_ (.A1(_1018_),
    .A2(_0409_),
    .B1(_1809_),
    .C1(_1810_),
    .D1(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__nand2_1 _5478_ (.A(_0430_),
    .B(_0731_),
    .Y(_1813_));
 sky130_fd_sc_hd__nand2_1 _5479_ (.A(_0434_),
    .B(_0733_),
    .Y(_1814_));
 sky130_fd_sc_hd__or2_1 _5480_ (.A(_0735_),
    .B(_0439_),
    .X(_1815_));
 sky130_fd_sc_hd__o2111a_1 _5481_ (.A1(_0365_),
    .A2(_0427_),
    .B1(_1813_),
    .C1(_1814_),
    .D1(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_0451_),
    .B(_0413_),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_0456_),
    .B(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .Y(_1818_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_1817_),
    .B(_1818_),
    .Y(_1819_));
 sky130_fd_sc_hd__a221oi_1 _5485_ (.A1(_1039_),
    .A2(_0445_),
    .B1(_0447_),
    .B2(_0461_),
    .C1(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__nand2_1 _5486_ (.A(_0471_),
    .B(_3168_),
    .Y(_1821_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(_0475_),
    .B(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_1822_));
 sky130_fd_sc_hd__nand2_1 _5488_ (.A(_1821_),
    .B(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__a221oi_1 _5489_ (.A1(_3171_),
    .A2(_0464_),
    .B1(_3174_),
    .B2(_0468_),
    .C1(_1823_),
    .Y(_1824_));
 sky130_fd_sc_hd__and4_1 _5490_ (.A(_1812_),
    .B(_1816_),
    .C(_1820_),
    .D(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__nand2_1 _5491_ (.A(_1808_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__nand2_1 _5492_ (.A(_0489_),
    .B(_0919_),
    .Y(_1827_));
 sky130_fd_sc_hd__o21ai_1 _5493_ (.A1(_0772_),
    .A2(_0486_),
    .B1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand2_1 _5494_ (.A(_0499_),
    .B(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_1829_));
 sky130_fd_sc_hd__nand2_1 _5495_ (.A(_0503_),
    .B(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _5496_ (.A(_1829_),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__a221oi_1 _5497_ (.A1(_0916_),
    .A2(_0494_),
    .B1(_0496_),
    .B2(_0518_),
    .C1(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5498_ (.A(_0509_),
    .B(_0538_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_0514_),
    .B(_0442_),
    .Y(_1834_));
 sky130_fd_sc_hd__and4b_1 _5500_ (.A_N(_1828_),
    .B(_1832_),
    .C(_1833_),
    .D(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__o22ai_1 _5501_ (.A1(_1202_),
    .A2(_0528_),
    .B1(_1334_),
    .B2(_0531_),
    .Y(_1836_));
 sky130_fd_sc_hd__a221oi_1 _5502_ (.A1(_0452_),
    .A2(_0521_),
    .B1(_0746_),
    .B2(_0525_),
    .C1(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__o22ai_1 _5503_ (.A1(_0437_),
    .A2(_0544_),
    .B1(_0743_),
    .B2(_0547_),
    .Y(_1838_));
 sky130_fd_sc_hd__a221oi_1 _5504_ (.A1(_0741_),
    .A2(_0537_),
    .B1(_0894_),
    .B2(_0541_),
    .C1(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__and3_1 _5505_ (.A(_1835_),
    .B(_1837_),
    .C(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__nand2_1 _5506_ (.A(_0563_),
    .B(_0573_),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _5507_ (.A(_0568_),
    .B(_0584_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _5508_ (.A(_1841_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__a221oi_1 _5509_ (.A1(_0577_),
    .A2(_0556_),
    .B1(_0781_),
    .B2(_0560_),
    .C1(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__nand2_1 _5510_ (.A(_0583_),
    .B(_0510_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2_1 _5511_ (.A(_0588_),
    .B(_1192_),
    .Y(_1846_));
 sky130_fd_sc_hd__nand2_1 _5512_ (.A(_1845_),
    .B(_1846_),
    .Y(_1847_));
 sky130_fd_sc_hd__a221oi_1 _5513_ (.A1(_0515_),
    .A2(_0576_),
    .B1(_0765_),
    .B2(_0580_),
    .C1(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _5514_ (.A(_0606_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_1849_));
 sky130_fd_sc_hd__o21ai_1 _5515_ (.A1(_0622_),
    .A2(_0603_),
    .B1(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__a221oi_1 _5516_ (.A1(_0615_),
    .A2(_0596_),
    .B1(_0589_),
    .B2(_0600_),
    .C1(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__inv_2 _5517_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_1852_));
 sky130_fd_sc_hd__o22ai_1 _5518_ (.A1(_1729_),
    .A2(_0621_),
    .B1(_1852_),
    .B2(_0624_),
    .Y(_1853_));
 sky130_fd_sc_hd__a221oi_1 _5519_ (.A1(_1210_),
    .A2(_0614_),
    .B1(_1055_),
    .B2(_0618_),
    .C1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__and4_1 _5520_ (.A(_1844_),
    .B(_1848_),
    .C(_1851_),
    .D(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__nand2_1 _5521_ (.A(_1840_),
    .B(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__nor2_1 _5522_ (.A(_1826_),
    .B(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(_0633_),
    .B(_0329_),
    .Y(_1858_));
 sky130_fd_sc_hd__nand3_2 _5524_ (.A(_1796_),
    .B(_1857_),
    .C(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__nor2_1 _5525_ (.A(_3212_),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__nor2_1 _5526_ (.A(_1738_),
    .B(_1860_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21ai_1 _5527_ (.A1(_3150_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .B1(_3161_),
    .Y(_1861_));
 sky130_fd_sc_hd__nand2_1 _5528_ (.A(_3236_),
    .B(_3255_),
    .Y(_1862_));
 sky130_fd_sc_hd__nand2_1 _5529_ (.A(_3244_),
    .B(_3250_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand2_1 _5530_ (.A(_1862_),
    .B(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__a221oi_1 _5531_ (.A1(_3432_),
    .A2(_3222_),
    .B1(_3439_),
    .B2(_3228_),
    .C1(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__nand2_1 _5532_ (.A(_3262_),
    .B(_3402_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _5533_ (.A(_3269_),
    .B(_3395_),
    .Y(_1867_));
 sky130_fd_sc_hd__nand2_1 _5534_ (.A(_1866_),
    .B(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__a221oi_1 _5535_ (.A1(_0675_),
    .A2(_3253_),
    .B1(_0836_),
    .B2(_3257_),
    .C1(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _5536_ (.A(_3294_),
    .B(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .Y(_1870_));
 sky130_fd_sc_hd__o21ai_1 _5537_ (.A1(_0964_),
    .A2(_3290_),
    .B1(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__a221oi_1 _5538_ (.A1(_3300_),
    .A2(_3280_),
    .B1(_3285_),
    .B2(_3306_),
    .C1(_1871_),
    .Y(_1872_));
 sky130_fd_sc_hd__o22ai_1 _5539_ (.A1(_3440_),
    .A2(_3313_),
    .B1(_0684_),
    .B2(_3317_),
    .Y(_1873_));
 sky130_fd_sc_hd__a221oi_1 _5540_ (.A1(_0991_),
    .A2(_3304_),
    .B1(_1130_),
    .B2(_3309_),
    .C1(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__and4_1 _5541_ (.A(_1865_),
    .B(_1869_),
    .C(_1872_),
    .D(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__nand2_1 _5542_ (.A(_3334_),
    .B(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_1876_));
 sky130_fd_sc_hd__o21ai_1 _5543_ (.A1(_0622_),
    .A2(_3122_),
    .B1(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__a221oi_1 _5544_ (.A1(_0551_),
    .A2(_3325_),
    .B1(_0557_),
    .B2(_3329_),
    .C1(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__nand2_1 _5545_ (.A(_3352_),
    .B(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .Y(_1879_));
 sky130_fd_sc_hd__o21ai_1 _5546_ (.A1(_0786_),
    .A2(_3349_),
    .B1(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__a221oi_1 _5547_ (.A1(_3336_),
    .A2(_3342_),
    .B1(_0657_),
    .B2(_3346_),
    .C1(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hd__nand2_1 _5548_ (.A(_3370_),
    .B(_3380_),
    .Y(_1882_));
 sky130_fd_sc_hd__o21ai_1 _5549_ (.A1(_0971_),
    .A2(_3367_),
    .B1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__a221oi_1 _5550_ (.A1(_3322_),
    .A2(_3360_),
    .B1(_3327_),
    .B2(_3364_),
    .C1(_1883_),
    .Y(_1884_));
 sky130_fd_sc_hd__nand2_1 _5551_ (.A(_3385_),
    .B(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_1885_));
 sky130_fd_sc_hd__nand2_1 _5552_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_1886_));
 sky130_fd_sc_hd__nand2_1 _5553_ (.A(_1885_),
    .B(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__a221oi_2 _5554_ (.A1(_0569_),
    .A2(_3378_),
    .B1(_0564_),
    .B2(_3382_),
    .C1(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__and4_1 _5555_ (.A(_1878_),
    .B(_1881_),
    .C(_1884_),
    .D(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__o22ai_1 _5556_ (.A1(_1767_),
    .A2(_3407_),
    .B1(_3422_),
    .B2(_3410_),
    .Y(_1890_));
 sky130_fd_sc_hd__a221oi_1 _5557_ (.A1(_0840_),
    .A2(_3400_),
    .B1(_3372_),
    .B2(_3404_),
    .C1(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__nand2_1 _5558_ (.A(_3426_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1892_));
 sky130_fd_sc_hd__o21ai_1 _5559_ (.A1(_0822_),
    .A2(_3423_),
    .B1(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__a221oi_1 _5560_ (.A1(_3354_),
    .A2(_3416_),
    .B1(_0662_),
    .B2(_3420_),
    .C1(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__nand2_1 _5561_ (.A(_3444_),
    .B(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .Y(_1895_));
 sky130_fd_sc_hd__o21ai_1 _5562_ (.A1(_1518_),
    .A2(_3441_),
    .B1(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__a221oi_1 _5563_ (.A1(_3449_),
    .A2(_3434_),
    .B1(_3437_),
    .B2(_3453_),
    .C1(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__nand2_1 _5564_ (.A(_3458_),
    .B(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_1898_));
 sky130_fd_sc_hd__nand2_1 _5565_ (.A(_3462_),
    .B(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .Y(_1899_));
 sky130_fd_sc_hd__nand2_1 _5566_ (.A(_1898_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__a221oi_1 _5567_ (.A1(_3340_),
    .A2(_3451_),
    .B1(_3344_),
    .B2(_3455_),
    .C1(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__and4_1 _5568_ (.A(_1891_),
    .B(_1894_),
    .C(_1897_),
    .D(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__nand2_1 _5569_ (.A(_3474_),
    .B(_3275_),
    .Y(_1903_));
 sky130_fd_sc_hd__nand2_1 _5570_ (.A(_3479_),
    .B(_3509_),
    .Y(_1904_));
 sky130_fd_sc_hd__or2_1 _5571_ (.A(_1146_),
    .B(_3484_),
    .X(_1905_));
 sky130_fd_sc_hd__o2111a_1 _5572_ (.A1(_0861_),
    .A2(_3471_),
    .B1(_1903_),
    .C1(_1904_),
    .D1(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__nand2_1 _5573_ (.A(_3495_),
    .B(_0865_),
    .Y(_1907_));
 sky130_fd_sc_hd__o221a_1 _5574_ (.A1(_3500_),
    .A2(_3489_),
    .B1(_1141_),
    .B2(_3492_),
    .C1(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__o22ai_1 _5575_ (.A1(_1100_),
    .A2(_3501_),
    .B1(_1237_),
    .B2(_3504_),
    .Y(_1909_));
 sky130_fd_sc_hd__a22o_1 _5576_ (.A1(_3507_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .B1(_3510_),
    .B2(_0801_),
    .X(_1910_));
 sky130_fd_sc_hd__nor2_1 _5577_ (.A(_1909_),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__nand2_1 _5578_ (.A(_0322_),
    .B(_3238_),
    .Y(_1912_));
 sky130_fd_sc_hd__nand2_1 _5579_ (.A(_0327_),
    .B(_3296_),
    .Y(_1913_));
 sky130_fd_sc_hd__nand2_1 _5580_ (.A(_0332_),
    .B(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _5581_ (.A(_0337_),
    .B(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .Y(_1915_));
 sky130_fd_sc_hd__and4_1 _5582_ (.A(_1912_),
    .B(_1913_),
    .C(_1914_),
    .D(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__and4_1 _5583_ (.A(_1906_),
    .B(_1908_),
    .C(_1911_),
    .D(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__and4_1 _5584_ (.A(_1875_),
    .B(_1889_),
    .C(_1902_),
    .D(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__nor2_1 _5585_ (.A(_0881_),
    .B(_0350_),
    .Y(_1919_));
 sky130_fd_sc_hd__a22o_1 _5586_ (.A1(_0353_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .B1(_0355_),
    .B2(_0796_),
    .X(_1920_));
 sky130_fd_sc_hd__a211oi_1 _5587_ (.A1(_3205_),
    .A2(_0347_),
    .B1(_1919_),
    .C1(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__nand2_1 _5588_ (.A(_0369_),
    .B(_3195_),
    .Y(_1922_));
 sky130_fd_sc_hd__o21ai_1 _5589_ (.A1(_1291_),
    .A2(_0366_),
    .B1(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__a221oi_1 _5590_ (.A1(_3199_),
    .A2(_0360_),
    .B1(_3202_),
    .B2(_0363_),
    .C1(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__o22ai_1 _5591_ (.A1(_0693_),
    .A2(_0381_),
    .B1(_3483_),
    .B2(_0384_),
    .Y(_1925_));
 sky130_fd_sc_hd__a221oi_1 _5592_ (.A1(_0339_),
    .A2(_0375_),
    .B1(_0329_),
    .B2(_0378_),
    .C1(_1925_),
    .Y(_1926_));
 sky130_fd_sc_hd__nand2_1 _5593_ (.A(_0398_),
    .B(_0701_),
    .Y(_1927_));
 sky130_fd_sc_hd__o21ai_1 _5594_ (.A1(_3468_),
    .A2(_0395_),
    .B1(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__a221oi_1 _5595_ (.A1(_0947_),
    .A2(_0389_),
    .B1(_3497_),
    .B2(_0392_),
    .C1(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__and4_1 _5596_ (.A(_1921_),
    .B(_1924_),
    .C(_1926_),
    .D(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__nand2_1 _5597_ (.A(_0411_),
    .B(_3180_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _5598_ (.A(_0416_),
    .B(_3186_),
    .Y(_1932_));
 sky130_fd_sc_hd__or2_1 _5599_ (.A(_0873_),
    .B(_0421_),
    .X(_1933_));
 sky130_fd_sc_hd__o2111a_1 _5600_ (.A1(_1157_),
    .A2(_0408_),
    .B1(_1931_),
    .C1(_1932_),
    .D1(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(_0429_),
    .B(_0418_),
    .Y(_1935_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_0433_),
    .B(_3152_),
    .Y(_1936_));
 sky130_fd_sc_hd__or2_1 _5603_ (.A(_0404_),
    .B(_0438_),
    .X(_1937_));
 sky130_fd_sc_hd__o2111a_1 _5604_ (.A1(_0720_),
    .A2(_0426_),
    .B1(_1935_),
    .C1(_1936_),
    .D1(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__nand2_1 _5605_ (.A(_0450_),
    .B(_0731_),
    .Y(_1939_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .Y(_1940_));
 sky130_fd_sc_hd__nand2_1 _5607_ (.A(_1939_),
    .B(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__a221oi_1 _5608_ (.A1(_0461_),
    .A2(_0444_),
    .B1(_0446_),
    .B2(_0465_),
    .C1(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5609_ (.A(_0470_),
    .B(_3171_),
    .Y(_1943_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(_0474_),
    .B(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_1944_));
 sky130_fd_sc_hd__nand2_1 _5611_ (.A(_1943_),
    .B(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__a221oi_1 _5612_ (.A1(_3174_),
    .A2(_0463_),
    .B1(_3177_),
    .B2(_0467_),
    .C1(_1945_),
    .Y(_1946_));
 sky130_fd_sc_hd__and4_1 _5613_ (.A(_1934_),
    .B(_1938_),
    .C(_1942_),
    .D(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__nand2_1 _5614_ (.A(_1930_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(_0488_),
    .B(_0534_),
    .Y(_1949_));
 sky130_fd_sc_hd__o21ai_1 _5616_ (.A1(_0923_),
    .A2(_0485_),
    .B1(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _5617_ (.A(_0498_),
    .B(_0919_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand2_1 _5618_ (.A(_0502_),
    .B(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_1952_));
 sky130_fd_sc_hd__nand2_1 _5619_ (.A(_1951_),
    .B(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__a221oi_1 _5620_ (.A1(_0518_),
    .A2(_0493_),
    .B1(_0495_),
    .B2(_0522_),
    .C1(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand2_1 _5621_ (.A(_0508_),
    .B(_0442_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand2_1 _5622_ (.A(_0513_),
    .B(_0448_),
    .Y(_1956_));
 sky130_fd_sc_hd__and4b_1 _5623_ (.A_N(_1950_),
    .B(_1954_),
    .C(_1955_),
    .D(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__o22ai_1 _5624_ (.A1(_1334_),
    .A2(_0527_),
    .B1(_1462_),
    .B2(_0530_),
    .Y(_1958_));
 sky130_fd_sc_hd__a221oi_1 _5625_ (.A1(_0746_),
    .A2(_0520_),
    .B1(_0739_),
    .B2(_0524_),
    .C1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__o22ai_1 _5626_ (.A1(_0743_),
    .A2(_0543_),
    .B1(_0425_),
    .B2(_0546_),
    .Y(_1960_));
 sky130_fd_sc_hd__a221oi_1 _5627_ (.A1(_0894_),
    .A2(_0536_),
    .B1(_1039_),
    .B2(_0540_),
    .C1(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__and3_1 _5628_ (.A(_1957_),
    .B(_1959_),
    .C(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__nand2_1 _5629_ (.A(_0562_),
    .B(_0577_),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_1 _5630_ (.A(_0567_),
    .B(_0573_),
    .Y(_1964_));
 sky130_fd_sc_hd__nand2_1 _5631_ (.A(_1963_),
    .B(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hd__a221oi_1 _5632_ (.A1(_0781_),
    .A2(_0555_),
    .B1(_0932_),
    .B2(_0559_),
    .C1(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_0582_),
    .B(_0515_),
    .Y(_1967_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(_0587_),
    .B(_0510_),
    .Y(_1968_));
 sky130_fd_sc_hd__nand2_1 _5635_ (.A(_1967_),
    .B(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__a221oi_1 _5636_ (.A1(_0765_),
    .A2(_0575_),
    .B1(_0916_),
    .B2(_0579_),
    .C1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _5637_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_1971_));
 sky130_fd_sc_hd__o21ai_1 _5638_ (.A1(_0790_),
    .A2(_0602_),
    .B1(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__a221oi_2 _5639_ (.A1(_0589_),
    .A2(_0595_),
    .B1(_0584_),
    .B2(_0599_),
    .C1(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__inv_2 _5640_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_1974_));
 sky130_fd_sc_hd__o22ai_1 _5641_ (.A1(_1852_),
    .A2(_0620_),
    .B1(_1974_),
    .B2(_0623_),
    .Y(_1975_));
 sky130_fd_sc_hd__a221oi_1 _5642_ (.A1(_1055_),
    .A2(_0613_),
    .B1(_1192_),
    .B2(_0617_),
    .C1(_1975_),
    .Y(_1976_));
 sky130_fd_sc_hd__and4_1 _5643_ (.A(_1966_),
    .B(_1970_),
    .C(_1973_),
    .D(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__nand2_1 _5644_ (.A(_1962_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__nor2_1 _5645_ (.A(_1948_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_0632_),
    .B(_0334_),
    .Y(_1980_));
 sky130_fd_sc_hd__nand3_1 _5647_ (.A(_1918_),
    .B(_1979_),
    .C(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__nor2_1 _5648_ (.A(_3149_),
    .B(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__nor2_1 _5649_ (.A(_1861_),
    .B(_1982_),
    .Y(_0287_));
 sky130_fd_sc_hd__o21ai_1 _5650_ (.A1(_3150_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .B1(_3161_),
    .Y(_1983_));
 sky130_fd_sc_hd__nand2_1 _5651_ (.A(_3236_),
    .B(_3432_),
    .Y(_1984_));
 sky130_fd_sc_hd__nand2_1 _5652_ (.A(_3244_),
    .B(_3255_),
    .Y(_1985_));
 sky130_fd_sc_hd__nand2_1 _5653_ (.A(_1984_),
    .B(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__a221oi_1 _5654_ (.A1(_3439_),
    .A2(_3222_),
    .B1(_0683_),
    .B2(_3228_),
    .C1(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__nand2_1 _5655_ (.A(_3262_),
    .B(_0675_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5656_ (.A(_3269_),
    .B(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _5657_ (.A(_1988_),
    .B(_1989_),
    .Y(_1990_));
 sky130_fd_sc_hd__a221oi_1 _5658_ (.A1(_0836_),
    .A2(_3253_),
    .B1(_3449_),
    .B2(_3257_),
    .C1(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand2_1 _5659_ (.A(_3294_),
    .B(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .Y(_1992_));
 sky130_fd_sc_hd__o21ai_1 _5660_ (.A1(_1104_),
    .A2(_3290_),
    .B1(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__a221oi_1 _5661_ (.A1(_3306_),
    .A2(_3280_),
    .B1(_3285_),
    .B2(_3271_),
    .C1(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__o22ai_1 _5662_ (.A1(_0684_),
    .A2(_3313_),
    .B1(_3406_),
    .B2(_3317_),
    .Y(_1995_));
 sky130_fd_sc_hd__a221oi_1 _5663_ (.A1(_1130_),
    .A2(_3304_),
    .B1(_3395_),
    .B2(_3309_),
    .C1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__and4_1 _5664_ (.A(_1987_),
    .B(_1991_),
    .C(_1994_),
    .D(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(_3334_),
    .B(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_1998_));
 sky130_fd_sc_hd__o21ai_1 _5666_ (.A1(_0790_),
    .A2(_3122_),
    .B1(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__a221oi_1 _5667_ (.A1(_0557_),
    .A2(_3325_),
    .B1(_0776_),
    .B2(_3329_),
    .C1(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__nand2_1 _5668_ (.A(_3352_),
    .B(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_2001_));
 sky130_fd_sc_hd__o21ai_1 _5669_ (.A1(_0937_),
    .A2(_3349_),
    .B1(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__a221oi_1 _5670_ (.A1(_0657_),
    .A2(_3342_),
    .B1(_0818_),
    .B2(_3346_),
    .C1(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_1 _5671_ (.A(_3370_),
    .B(_3322_),
    .Y(_2004_));
 sky130_fd_sc_hd__o21ai_1 _5672_ (.A1(_1111_),
    .A2(_3367_),
    .B1(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__a221oi_1 _5673_ (.A1(_3327_),
    .A2(_3360_),
    .B1(_3336_),
    .B2(_3364_),
    .C1(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__nand2_1 _5674_ (.A(_3385_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_2007_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_2008_));
 sky130_fd_sc_hd__nand2_1 _5676_ (.A(_2007_),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__a221oi_1 _5677_ (.A1(_0564_),
    .A2(_3378_),
    .B1(_0551_),
    .B2(_3382_),
    .C1(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__and4_1 _5678_ (.A(_2000_),
    .B(_2003_),
    .C(_2006_),
    .D(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__o22ai_1 _5679_ (.A1(_3422_),
    .A2(_3407_),
    .B1(_3366_),
    .B2(_3410_),
    .Y(_2012_));
 sky130_fd_sc_hd__a221oi_1 _5680_ (.A1(_3372_),
    .A2(_3400_),
    .B1(_3358_),
    .B2(_3404_),
    .C1(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hd__nand2_1 _5681_ (.A(_3426_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_2014_));
 sky130_fd_sc_hd__o21ai_1 _5682_ (.A1(_0971_),
    .A2(_3423_),
    .B1(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__a221oi_1 _5683_ (.A1(_0662_),
    .A2(_3416_),
    .B1(_0823_),
    .B2(_3420_),
    .C1(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _5684_ (.A(_3444_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_2017_));
 sky130_fd_sc_hd__o21ai_1 _5685_ (.A1(_1644_),
    .A2(_3441_),
    .B1(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__a221oi_1 _5686_ (.A1(_3453_),
    .A2(_3434_),
    .B1(_3437_),
    .B2(_3414_),
    .C1(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _5687_ (.A(_3458_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_2020_));
 sky130_fd_sc_hd__nand2_1 _5688_ (.A(_3462_),
    .B(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_1 _5689_ (.A(_2020_),
    .B(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__a221oi_1 _5690_ (.A1(_3344_),
    .A2(_3451_),
    .B1(_3354_),
    .B2(_3455_),
    .C1(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__and4_1 _5691_ (.A(_2013_),
    .B(_2016_),
    .C(_2019_),
    .D(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__nand2_1 _5692_ (.A(_3474_),
    .B(_3287_),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _5693_ (.A(_3479_),
    .B(_3512_),
    .Y(_2026_));
 sky130_fd_sc_hd__or2_1 _5694_ (.A(_3288_),
    .B(_3484_),
    .X(_2027_));
 sky130_fd_sc_hd__o2111a_1 _5695_ (.A1(_1007_),
    .A2(_3471_),
    .B1(_2025_),
    .C1(_2026_),
    .D1(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__nand2_1 _5696_ (.A(_3495_),
    .B(_3509_),
    .Y(_2029_));
 sky130_fd_sc_hd__o221a_1 _5697_ (.A1(_3503_),
    .A2(_3489_),
    .B1(_3500_),
    .B2(_3492_),
    .C1(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__o22ai_1 _5698_ (.A1(_1237_),
    .A2(_3501_),
    .B1(_3311_),
    .B2(_3504_),
    .Y(_2031_));
 sky130_fd_sc_hd__a22o_1 _5699_ (.A1(_3507_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .B1(_3510_),
    .B2(_3300_),
    .X(_2032_));
 sky130_fd_sc_hd__nor2_1 _5700_ (.A(_2031_),
    .B(_2032_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand2_1 _5701_ (.A(_0322_),
    .B(_3213_),
    .Y(_2034_));
 sky130_fd_sc_hd__nand2_1 _5702_ (.A(_0327_),
    .B(_3246_),
    .Y(_2035_));
 sky130_fd_sc_hd__nand2_1 _5703_ (.A(_0332_),
    .B(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .Y(_2036_));
 sky130_fd_sc_hd__nand2_1 _5704_ (.A(_0337_),
    .B(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .Y(_2037_));
 sky130_fd_sc_hd__and4_1 _5705_ (.A(_2034_),
    .B(_2035_),
    .C(_2036_),
    .D(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__and4_1 _5706_ (.A(_2028_),
    .B(_2030_),
    .C(_2033_),
    .D(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__and4_1 _5707_ (.A(_1997_),
    .B(_2011_),
    .C(_2024_),
    .D(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__nor2_1 _5708_ (.A(_1026_),
    .B(_0350_),
    .Y(_2041_));
 sky130_fd_sc_hd__a22o_1 _5709_ (.A1(_0353_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .B1(_0355_),
    .B2(_0947_),
    .X(_2042_));
 sky130_fd_sc_hd__a211oi_1 _5710_ (.A1(_3208_),
    .A2(_0347_),
    .B1(_2041_),
    .C1(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_0369_),
    .B(_3199_),
    .Y(_2044_));
 sky130_fd_sc_hd__o21ai_1 _5712_ (.A1(_0394_),
    .A2(_0366_),
    .B1(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__a221oi_1 _5713_ (.A1(_3202_),
    .A2(_0360_),
    .B1(_3205_),
    .B2(_0363_),
    .C1(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__o22ai_1 _5714_ (.A1(_3483_),
    .A2(_0381_),
    .B1(_0697_),
    .B2(_0384_),
    .Y(_2047_));
 sky130_fd_sc_hd__a221oi_1 _5715_ (.A1(_0329_),
    .A2(_0375_),
    .B1(_0334_),
    .B2(_0378_),
    .C1(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__nand2_1 _5716_ (.A(_0398_),
    .B(_0695_),
    .Y(_2049_));
 sky130_fd_sc_hd__o21ai_1 _5717_ (.A1(_0693_),
    .A2(_0395_),
    .B1(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__a221oi_1 _5718_ (.A1(_3497_),
    .A2(_0389_),
    .B1(_0701_),
    .B2(_0392_),
    .C1(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__and4_1 _5719_ (.A(_2043_),
    .B(_2046_),
    .C(_2048_),
    .D(_2051_),
    .X(_2052_));
 sky130_fd_sc_hd__nand2_1 _5720_ (.A(_0411_),
    .B(_3183_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _5721_ (.A(_0416_),
    .B(_3189_),
    .Y(_2054_));
 sky130_fd_sc_hd__or2_1 _5722_ (.A(_1018_),
    .B(_0421_),
    .X(_2055_));
 sky130_fd_sc_hd__o2111a_1 _5723_ (.A1(_1291_),
    .A2(_0408_),
    .B1(_2053_),
    .C1(_2054_),
    .D1(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__nand2_1 _5724_ (.A(_0429_),
    .B(_0733_),
    .Y(_2057_));
 sky130_fd_sc_hd__nand2_1 _5725_ (.A(_0433_),
    .B(_3163_),
    .Y(_2058_));
 sky130_fd_sc_hd__or2_1 _5726_ (.A(_0365_),
    .B(_0438_),
    .X(_2059_));
 sky130_fd_sc_hd__o2111a_1 _5727_ (.A1(_0877_),
    .A2(_0426_),
    .B1(_2057_),
    .C1(_2058_),
    .D1(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__nand2_1 _5728_ (.A(_0450_),
    .B(_0418_),
    .Y(_2061_));
 sky130_fd_sc_hd__nand2_1 _5729_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .Y(_2062_));
 sky130_fd_sc_hd__nand2_1 _5730_ (.A(_2061_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__a221oi_1 _5731_ (.A1(_0465_),
    .A2(_0444_),
    .B1(_0446_),
    .B2(_0413_),
    .C1(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__nand2_1 _5732_ (.A(_0470_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_2065_));
 sky130_fd_sc_hd__nand2_1 _5733_ (.A(_0474_),
    .B(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_2066_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_2065_),
    .B(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__a221oi_1 _5735_ (.A1(_3177_),
    .A2(_0463_),
    .B1(_3180_),
    .B2(_0467_),
    .C1(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__and4_1 _5736_ (.A(_2056_),
    .B(_2060_),
    .C(_2064_),
    .D(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__nand2_1 _5737_ (.A(_2052_),
    .B(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__nand2_1 _5738_ (.A(_0488_),
    .B(_0538_),
    .Y(_2071_));
 sky130_fd_sc_hd__o21ai_1 _5739_ (.A1(_1065_),
    .A2(_0485_),
    .B1(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__nand2_1 _5740_ (.A(_0498_),
    .B(_0534_),
    .Y(_2073_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(_0502_),
    .B(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_2074_));
 sky130_fd_sc_hd__nand2_1 _5742_ (.A(_2073_),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__a221oi_1 _5743_ (.A1(_0522_),
    .A2(_0493_),
    .B1(_0495_),
    .B2(_0768_),
    .C1(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand2_1 _5744_ (.A(_0508_),
    .B(_0448_),
    .Y(_2077_));
 sky130_fd_sc_hd__nand2_1 _5745_ (.A(_0513_),
    .B(_0457_),
    .Y(_2078_));
 sky130_fd_sc_hd__and4b_1 _5746_ (.A_N(_2072_),
    .B(_2076_),
    .C(_2077_),
    .D(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__o22ai_1 _5747_ (.A1(_1462_),
    .A2(_0527_),
    .B1(_1589_),
    .B2(_0530_),
    .Y(_2080_));
 sky130_fd_sc_hd__a221oi_1 _5748_ (.A1(_0739_),
    .A2(_0520_),
    .B1(_0435_),
    .B2(_0524_),
    .C1(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__o22ai_1 _5749_ (.A1(_0425_),
    .A2(_0543_),
    .B1(_0738_),
    .B2(_0546_),
    .Y(_2082_));
 sky130_fd_sc_hd__a221oi_1 _5750_ (.A1(_1039_),
    .A2(_0536_),
    .B1(_0461_),
    .B2(_0540_),
    .C1(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__and3_1 _5751_ (.A(_2079_),
    .B(_2081_),
    .C(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__nand2_1 _5752_ (.A(_0562_),
    .B(_0781_),
    .Y(_2085_));
 sky130_fd_sc_hd__nand2_1 _5753_ (.A(_0567_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_2086_));
 sky130_fd_sc_hd__nand2_1 _5754_ (.A(_2085_),
    .B(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__a221oi_1 _5755_ (.A1(_0932_),
    .A2(_0555_),
    .B1(_1073_),
    .B2(_0559_),
    .C1(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2_1 _5756_ (.A(_0582_),
    .B(_0765_),
    .Y(_2089_));
 sky130_fd_sc_hd__nand2_1 _5757_ (.A(_0587_),
    .B(_0515_),
    .Y(_2090_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(_2089_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__a221oi_1 _5759_ (.A1(_0916_),
    .A2(_0575_),
    .B1(_0518_),
    .B2(_0579_),
    .C1(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_2093_));
 sky130_fd_sc_hd__o21ai_1 _5761_ (.A1(_0941_),
    .A2(_0602_),
    .B1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__a221oi_2 _5762_ (.A1(_0584_),
    .A2(_0595_),
    .B1(_0573_),
    .B2(_0599_),
    .C1(_2094_),
    .Y(_2095_));
 sky130_fd_sc_hd__inv_2 _5763_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_2096_));
 sky130_fd_sc_hd__o22ai_1 _5764_ (.A1(_1974_),
    .A2(_0620_),
    .B1(_2096_),
    .B2(_0623_),
    .Y(_2097_));
 sky130_fd_sc_hd__a221oi_1 _5765_ (.A1(_1192_),
    .A2(_0613_),
    .B1(_0510_),
    .B2(_0617_),
    .C1(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__and4_1 _5766_ (.A(_2088_),
    .B(_2092_),
    .C(_2095_),
    .D(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(_2084_),
    .B(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__nor2_1 _5768_ (.A(_2070_),
    .B(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__nand2_1 _5769_ (.A(_0632_),
    .B(_0324_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand3_1 _5770_ (.A(_2040_),
    .B(_2101_),
    .C(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__nor2_1 _5771_ (.A(_3149_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__nor2_1 _5772_ (.A(_1983_),
    .B(_2104_),
    .Y(_0286_));
 sky130_fd_sc_hd__o21ai_1 _5773_ (.A1(_3150_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .B1(_3161_),
    .Y(_2105_));
 sky130_fd_sc_hd__nand2_1 _5774_ (.A(_3236_),
    .B(_3439_),
    .Y(_2106_));
 sky130_fd_sc_hd__nand2_1 _5775_ (.A(_3244_),
    .B(_3432_),
    .Y(_2107_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(_2106_),
    .B(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__a221oi_1 _5777_ (.A1(_0683_),
    .A2(_3222_),
    .B1(_0844_),
    .B2(_3228_),
    .C1(_2108_),
    .Y(_2109_));
 sky130_fd_sc_hd__nand2_1 _5778_ (.A(_3262_),
    .B(_0836_),
    .Y(_2110_));
 sky130_fd_sc_hd__nand2_1 _5779_ (.A(_3269_),
    .B(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_1 _5780_ (.A(_2110_),
    .B(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__a221oi_1 _5781_ (.A1(_3449_),
    .A2(_3253_),
    .B1(_3453_),
    .B2(_3257_),
    .C1(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__nand2_1 _5782_ (.A(_3294_),
    .B(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .Y(_2114_));
 sky130_fd_sc_hd__o21ai_1 _5783_ (.A1(_1241_),
    .A2(_3290_),
    .B1(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__a221oi_1 _5784_ (.A1(_3271_),
    .A2(_3280_),
    .B1(_3285_),
    .B2(_3264_),
    .C1(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__o22ai_1 _5785_ (.A1(_3406_),
    .A2(_3313_),
    .B1(_3409_),
    .B2(_3317_),
    .Y(_2117_));
 sky130_fd_sc_hd__a221oi_1 _5786_ (.A1(_3395_),
    .A2(_3304_),
    .B1(_3402_),
    .B2(_3309_),
    .C1(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__and4_1 _5787_ (.A(_2109_),
    .B(_2113_),
    .C(_2116_),
    .D(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__nand2_1 _5788_ (.A(_3334_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_2120_));
 sky130_fd_sc_hd__o21ai_1 _5789_ (.A1(_0941_),
    .A2(_3122_),
    .B1(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__a221oi_1 _5790_ (.A1(_0776_),
    .A2(_3325_),
    .B1(_0927_),
    .B2(_3329_),
    .C1(_2121_),
    .Y(_2122_));
 sky130_fd_sc_hd__nand2_1 _5791_ (.A(_3352_),
    .B(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_2123_));
 sky130_fd_sc_hd__o21ai_1 _5792_ (.A1(_1078_),
    .A2(_3349_),
    .B1(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__a221oi_1 _5793_ (.A1(_0818_),
    .A2(_3342_),
    .B1(_0607_),
    .B2(_3346_),
    .C1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__nand2_1 _5794_ (.A(_3370_),
    .B(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .Y(_2126_));
 sky130_fd_sc_hd__o21ai_1 _5795_ (.A1(_1248_),
    .A2(_3367_),
    .B1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__a221oi_1 _5796_ (.A1(_3336_),
    .A2(_3360_),
    .B1(_0657_),
    .B2(_3364_),
    .C1(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__nand2_1 _5797_ (.A(_3385_),
    .B(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_2129_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_2130_));
 sky130_fd_sc_hd__nand2_1 _5799_ (.A(_2129_),
    .B(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__a221oi_1 _5800_ (.A1(_0551_),
    .A2(_3378_),
    .B1(_0557_),
    .B2(_3382_),
    .C1(_2131_),
    .Y(_2132_));
 sky130_fd_sc_hd__and4_1 _5801_ (.A(_2122_),
    .B(_2125_),
    .C(_2128_),
    .D(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__o22ai_1 _5802_ (.A1(_3366_),
    .A2(_3407_),
    .B1(_0666_),
    .B2(_3410_),
    .Y(_2134_));
 sky130_fd_sc_hd__a221oi_1 _5803_ (.A1(_3358_),
    .A2(_3400_),
    .B1(_3362_),
    .B2(_3404_),
    .C1(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__nand2_1 _5804_ (.A(_3426_),
    .B(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .Y(_2136_));
 sky130_fd_sc_hd__o21ai_1 _5805_ (.A1(_1111_),
    .A2(_3423_),
    .B1(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__a221oi_1 _5806_ (.A1(_0823_),
    .A2(_3416_),
    .B1(_0972_),
    .B2(_3420_),
    .C1(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__nand2_1 _5807_ (.A(_3444_),
    .B(_0679_),
    .Y(_2139_));
 sky130_fd_sc_hd__o21ai_1 _5808_ (.A1(_1767_),
    .A2(_3441_),
    .B1(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__a221oi_1 _5809_ (.A1(_3414_),
    .A2(_3434_),
    .B1(_3437_),
    .B2(_3418_),
    .C1(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(_3458_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_2142_));
 sky130_fd_sc_hd__nand2_1 _5811_ (.A(_3462_),
    .B(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .Y(_2143_));
 sky130_fd_sc_hd__nand2_1 _5812_ (.A(_2142_),
    .B(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__a221oi_1 _5813_ (.A1(_3354_),
    .A2(_3451_),
    .B1(_0662_),
    .B2(_3455_),
    .C1(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__and4_1 _5814_ (.A(_2135_),
    .B(_2138_),
    .C(_2141_),
    .D(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(_3474_),
    .B(_0648_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand2_1 _5816_ (.A(_3479_),
    .B(_3275_),
    .Y(_2148_));
 sky130_fd_sc_hd__or2_1 _5817_ (.A(_0649_),
    .B(_3484_),
    .X(_2149_));
 sky130_fd_sc_hd__o2111a_1 _5818_ (.A1(_1146_),
    .A2(_3471_),
    .B1(_2147_),
    .C1(_2148_),
    .D1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_3495_),
    .B(_3512_),
    .Y(_2151_));
 sky130_fd_sc_hd__o221a_1 _5820_ (.A1(_0704_),
    .A2(_3489_),
    .B1(_3503_),
    .B2(_3492_),
    .C1(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__o22ai_1 _5821_ (.A1(_3311_),
    .A2(_3501_),
    .B1(_3315_),
    .B2(_3504_),
    .Y(_2153_));
 sky130_fd_sc_hd__a22o_1 _5822_ (.A1(_3507_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .B1(_3510_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .X(_2154_));
 sky130_fd_sc_hd__nor2_1 _5823_ (.A(_2153_),
    .B(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_0322_),
    .B(_3224_),
    .Y(_2156_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_0327_),
    .B(_3238_),
    .Y(_2157_));
 sky130_fd_sc_hd__nand2_1 _5826_ (.A(_0332_),
    .B(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .Y(_2158_));
 sky130_fd_sc_hd__nand2_1 _5827_ (.A(_0337_),
    .B(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .Y(_2159_));
 sky130_fd_sc_hd__and4_1 _5828_ (.A(_2156_),
    .B(_2157_),
    .C(_2158_),
    .D(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__and4_1 _5829_ (.A(_2150_),
    .B(_2152_),
    .C(_2155_),
    .D(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__and4_1 _5830_ (.A(_2119_),
    .B(_2133_),
    .C(_2146_),
    .D(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__nor2_1 _5831_ (.A(_3491_),
    .B(_0350_),
    .Y(_2163_));
 sky130_fd_sc_hd__a22o_1 _5832_ (.A1(_0353_),
    .A2(_0947_),
    .B1(_0355_),
    .B2(_3497_),
    .X(_2164_));
 sky130_fd_sc_hd__a211oi_1 _5833_ (.A1(_0634_),
    .A2(_0347_),
    .B1(_2163_),
    .C1(_2164_),
    .Y(_2165_));
 sky130_fd_sc_hd__nand2_1 _5834_ (.A(_0369_),
    .B(_3202_),
    .Y(_2166_));
 sky130_fd_sc_hd__o21ai_1 _5835_ (.A1(_0380_),
    .A2(_0366_),
    .B1(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__a221oi_1 _5836_ (.A1(_3205_),
    .A2(_0360_),
    .B1(_3208_),
    .B2(_0363_),
    .C1(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__o22ai_1 _5837_ (.A1(_0697_),
    .A2(_0381_),
    .B1(_0855_),
    .B2(_0384_),
    .Y(_2169_));
 sky130_fd_sc_hd__a221oi_1 _5838_ (.A1(_0334_),
    .A2(_0375_),
    .B1(_0324_),
    .B2(_0378_),
    .C1(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__nand2_1 _5839_ (.A(_0398_),
    .B(_3476_),
    .Y(_2171_));
 sky130_fd_sc_hd__o21ai_1 _5840_ (.A1(_3483_),
    .A2(_0395_),
    .B1(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__a221oi_1 _5841_ (.A1(_0701_),
    .A2(_0389_),
    .B1(_0695_),
    .B2(_0392_),
    .C1(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__and4_1 _5842_ (.A(_2165_),
    .B(_2168_),
    .C(_2170_),
    .D(_2173_),
    .X(_2174_));
 sky130_fd_sc_hd__nand2_1 _5843_ (.A(_0411_),
    .B(_3186_),
    .Y(_2175_));
 sky130_fd_sc_hd__nand2_1 _5844_ (.A(_0416_),
    .B(_3192_),
    .Y(_2176_));
 sky130_fd_sc_hd__or2_1 _5845_ (.A(_1157_),
    .B(_0421_),
    .X(_2177_));
 sky130_fd_sc_hd__o2111a_1 _5846_ (.A1(_0394_),
    .A2(_0408_),
    .B1(_2175_),
    .C1(_2176_),
    .D1(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_0429_),
    .B(_3152_),
    .Y(_2179_));
 sky130_fd_sc_hd__nand2_1 _5848_ (.A(_0433_),
    .B(_3168_),
    .Y(_2180_));
 sky130_fd_sc_hd__or2_1 _5849_ (.A(_0720_),
    .B(_0438_),
    .X(_2181_));
 sky130_fd_sc_hd__o2111a_1 _5850_ (.A1(_1022_),
    .A2(_0426_),
    .B1(_2179_),
    .C1(_2180_),
    .D1(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__nand2_1 _5851_ (.A(_0450_),
    .B(_0733_),
    .Y(_2183_));
 sky130_fd_sc_hd__nand2_1 _5852_ (.A(_0455_),
    .B(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .Y(_2184_));
 sky130_fd_sc_hd__nand2_1 _5853_ (.A(_2183_),
    .B(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__a221oi_1 _5854_ (.A1(_0413_),
    .A2(_0444_),
    .B1(_0446_),
    .B2(_0731_),
    .C1(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_0470_),
    .B(_3177_),
    .Y(_2187_));
 sky130_fd_sc_hd__nand2_1 _5856_ (.A(_0474_),
    .B(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_2188_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(_2187_),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__a221oi_1 _5858_ (.A1(_3180_),
    .A2(_0463_),
    .B1(_3183_),
    .B2(_0467_),
    .C1(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__and4_1 _5859_ (.A(_2178_),
    .B(_2182_),
    .C(_2186_),
    .D(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__nand2_1 _5860_ (.A(_2174_),
    .B(_2191_),
    .Y(_2192_));
 sky130_fd_sc_hd__nand2_1 _5861_ (.A(_0488_),
    .B(_0442_),
    .Y(_2193_));
 sky130_fd_sc_hd__o21ai_1 _5862_ (.A1(_1202_),
    .A2(_0485_),
    .B1(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__nand2_1 _5863_ (.A(_0498_),
    .B(_0538_),
    .Y(_2195_));
 sky130_fd_sc_hd__nand2_1 _5864_ (.A(_0502_),
    .B(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_2196_));
 sky130_fd_sc_hd__nand2_1 _5865_ (.A(_2195_),
    .B(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__a221oi_1 _5866_ (.A1(_0768_),
    .A2(_0493_),
    .B1(_0495_),
    .B2(_0919_),
    .C1(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__nand2_1 _5867_ (.A(_0508_),
    .B(_0457_),
    .Y(_2199_));
 sky130_fd_sc_hd__nand2_1 _5868_ (.A(_0513_),
    .B(_0452_),
    .Y(_2200_));
 sky130_fd_sc_hd__and4b_1 _5869_ (.A_N(_2194_),
    .B(_2198_),
    .C(_2199_),
    .D(_2200_),
    .X(_2201_));
 sky130_fd_sc_hd__o22ai_1 _5870_ (.A1(_1589_),
    .A2(_0527_),
    .B1(_0437_),
    .B2(_0530_),
    .Y(_2202_));
 sky130_fd_sc_hd__a221oi_1 _5871_ (.A1(_0435_),
    .A2(_0520_),
    .B1(_0741_),
    .B2(_0524_),
    .C1(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__o22ai_1 _5872_ (.A1(_0738_),
    .A2(_0543_),
    .B1(_0892_),
    .B2(_0546_),
    .Y(_2204_));
 sky130_fd_sc_hd__a221oi_1 _5873_ (.A1(_0461_),
    .A2(_0536_),
    .B1(_0465_),
    .B2(_0540_),
    .C1(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__and3_1 _5874_ (.A(_2201_),
    .B(_2203_),
    .C(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__nand2_1 _5875_ (.A(_0562_),
    .B(_0932_),
    .Y(_2207_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_0567_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_2208_));
 sky130_fd_sc_hd__nand2_1 _5877_ (.A(_2207_),
    .B(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hd__a221oi_1 _5878_ (.A1(_1073_),
    .A2(_0555_),
    .B1(_1210_),
    .B2(_0559_),
    .C1(_2209_),
    .Y(_2210_));
 sky130_fd_sc_hd__nand2_1 _5879_ (.A(_0582_),
    .B(_0916_),
    .Y(_2211_));
 sky130_fd_sc_hd__nand2_1 _5880_ (.A(_0587_),
    .B(_0765_),
    .Y(_2212_));
 sky130_fd_sc_hd__nand2_1 _5881_ (.A(_2211_),
    .B(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__a221oi_1 _5882_ (.A1(_0518_),
    .A2(_0575_),
    .B1(_0522_),
    .B2(_0579_),
    .C1(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__nand2_1 _5883_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_2215_));
 sky130_fd_sc_hd__o21ai_1 _5884_ (.A1(_1082_),
    .A2(_0602_),
    .B1(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__a221oi_1 _5885_ (.A1(_0573_),
    .A2(_0595_),
    .B1(_0577_),
    .B2(_0599_),
    .C1(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__o22ai_1 _5886_ (.A1(_2096_),
    .A2(_0620_),
    .B1(_0481_),
    .B2(_0623_),
    .Y(_2218_));
 sky130_fd_sc_hd__a221oi_1 _5887_ (.A1(_0510_),
    .A2(_0613_),
    .B1(_0515_),
    .B2(_0617_),
    .C1(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__and4_1 _5888_ (.A(_2210_),
    .B(_2214_),
    .C(_2217_),
    .D(_2219_),
    .X(_2220_));
 sky130_fd_sc_hd__nand2_1 _5889_ (.A(_2206_),
    .B(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hd__nor2_1 _5890_ (.A(_2192_),
    .B(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__nand2_1 _5891_ (.A(_0632_),
    .B(_0708_),
    .Y(_2223_));
 sky130_fd_sc_hd__nand3_1 _5892_ (.A(_2162_),
    .B(_2222_),
    .C(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__nor2_1 _5893_ (.A(_3149_),
    .B(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__nor2_1 _5894_ (.A(_2105_),
    .B(_2225_),
    .Y(_0285_));
 sky130_fd_sc_hd__o21ai_1 _5895_ (.A1(_3150_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_3161_),
    .Y(_2226_));
 sky130_fd_sc_hd__nand2_1 _5896_ (.A(_3236_),
    .B(_0683_),
    .Y(_2227_));
 sky130_fd_sc_hd__nand2_1 _5897_ (.A(_3244_),
    .B(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_2228_));
 sky130_fd_sc_hd__nand2_1 _5898_ (.A(_2227_),
    .B(_2228_),
    .Y(_2229_));
 sky130_fd_sc_hd__a221oi_1 _5899_ (.A1(_0844_),
    .A2(_3222_),
    .B1(_0991_),
    .B2(_3228_),
    .C1(_2229_),
    .Y(_2230_));
 sky130_fd_sc_hd__nand2_1 _5900_ (.A(_3262_),
    .B(_3449_),
    .Y(_2231_));
 sky130_fd_sc_hd__nand2_1 _5901_ (.A(_3269_),
    .B(_0836_),
    .Y(_2232_));
 sky130_fd_sc_hd__nand2_1 _5902_ (.A(_2231_),
    .B(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__a221oi_1 _5903_ (.A1(_3453_),
    .A2(_3253_),
    .B1(_3414_),
    .B2(_3257_),
    .C1(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__nand2_1 _5904_ (.A(_3294_),
    .B(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .Y(_2235_));
 sky130_fd_sc_hd__o21ai_1 _5905_ (.A1(_1371_),
    .A2(_3290_),
    .B1(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__a221oi_1 _5906_ (.A1(_3264_),
    .A2(_3280_),
    .B1(_3285_),
    .B2(_3250_),
    .C1(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__o22ai_1 _5907_ (.A1(_3409_),
    .A2(_3313_),
    .B1(_0676_),
    .B2(_3317_),
    .Y(_2238_));
 sky130_fd_sc_hd__a221oi_1 _5908_ (.A1(_3402_),
    .A2(_3304_),
    .B1(_0675_),
    .B2(_3309_),
    .C1(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__and4_1 _5909_ (.A(_2230_),
    .B(_2234_),
    .C(_2237_),
    .D(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__nand2_1 _5910_ (.A(_3334_),
    .B(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_2241_));
 sky130_fd_sc_hd__o21ai_1 _5911_ (.A1(_1082_),
    .A2(_3122_),
    .B1(_2241_),
    .Y(_2242_));
 sky130_fd_sc_hd__a221oi_1 _5912_ (.A1(_0927_),
    .A2(_3325_),
    .B1(_0611_),
    .B2(_3329_),
    .C1(_2242_),
    .Y(_2243_));
 sky130_fd_sc_hd__nand2_1 _5913_ (.A(_3352_),
    .B(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_2244_));
 sky130_fd_sc_hd__o21ai_1 _5914_ (.A1(_1215_),
    .A2(_3349_),
    .B1(_2244_),
    .Y(_2245_));
 sky130_fd_sc_hd__a221oi_1 _5915_ (.A1(_0607_),
    .A2(_3342_),
    .B1(_0593_),
    .B2(_3346_),
    .C1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__nand2_1 _5916_ (.A(_3370_),
    .B(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .Y(_2247_));
 sky130_fd_sc_hd__o21ai_1 _5917_ (.A1(_1378_),
    .A2(_3367_),
    .B1(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__a221oi_1 _5918_ (.A1(_0657_),
    .A2(_3360_),
    .B1(_0818_),
    .B2(_3364_),
    .C1(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_3385_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_2250_));
 sky130_fd_sc_hd__nand2_1 _5920_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_2251_));
 sky130_fd_sc_hd__nand2_1 _5921_ (.A(_2250_),
    .B(_2251_),
    .Y(_2252_));
 sky130_fd_sc_hd__a221oi_2 _5922_ (.A1(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .A2(_3378_),
    .B1(_0776_),
    .B2(_3382_),
    .C1(_2252_),
    .Y(_2253_));
 sky130_fd_sc_hd__and4_1 _5923_ (.A(_2243_),
    .B(_2246_),
    .C(_2249_),
    .D(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__o22ai_1 _5924_ (.A1(_0666_),
    .A2(_3407_),
    .B1(_0827_),
    .B2(_3410_),
    .Y(_2255_));
 sky130_fd_sc_hd__a221oi_1 _5925_ (.A1(_3362_),
    .A2(_3400_),
    .B1(_3340_),
    .B2(_3404_),
    .C1(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__nand2_1 _5926_ (.A(_3426_),
    .B(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .Y(_2257_));
 sky130_fd_sc_hd__o21ai_1 _5927_ (.A1(_1248_),
    .A2(_3423_),
    .B1(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__a221oi_1 _5928_ (.A1(_0972_),
    .A2(_3416_),
    .B1(_3376_),
    .B2(_3420_),
    .C1(_2258_),
    .Y(_2259_));
 sky130_fd_sc_hd__nand2_1 _5929_ (.A(_3444_),
    .B(_0840_),
    .Y(_2260_));
 sky130_fd_sc_hd__o21ai_1 _5930_ (.A1(_3422_),
    .A2(_3441_),
    .B1(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__a221oi_1 _5931_ (.A1(_3418_),
    .A2(_3434_),
    .B1(_3437_),
    .B2(_3428_),
    .C1(_2261_),
    .Y(_2262_));
 sky130_fd_sc_hd__nand2_1 _5932_ (.A(_3458_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_2263_));
 sky130_fd_sc_hd__nand2_1 _5933_ (.A(_3462_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_2264_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(_2263_),
    .B(_2264_),
    .Y(_2265_));
 sky130_fd_sc_hd__a221oi_1 _5935_ (.A1(_0662_),
    .A2(_3451_),
    .B1(_0823_),
    .B2(_3455_),
    .C1(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__and4_1 _5936_ (.A(_2256_),
    .B(_2259_),
    .C(_2262_),
    .D(_2266_),
    .X(_2267_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(_3474_),
    .B(_3296_),
    .Y(_2268_));
 sky130_fd_sc_hd__nand2_1 _5938_ (.A(_3479_),
    .B(_3287_),
    .Y(_2269_));
 sky130_fd_sc_hd__or2_1 _5939_ (.A(_0810_),
    .B(_3484_),
    .X(_2270_));
 sky130_fd_sc_hd__o2111a_1 _5940_ (.A1(_3288_),
    .A2(_3471_),
    .B1(_2268_),
    .C1(_2269_),
    .D1(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__nand2_1 _5941_ (.A(_3495_),
    .B(_3275_),
    .Y(_2272_));
 sky130_fd_sc_hd__o221a_1 _5942_ (.A1(_0861_),
    .A2(_3489_),
    .B1(_0704_),
    .B2(_3492_),
    .C1(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__o22ai_1 _5943_ (.A1(_3315_),
    .A2(_3501_),
    .B1(_0653_),
    .B2(_3504_),
    .Y(_2274_));
 sky130_fd_sc_hd__a22o_1 _5944_ (.A1(_3507_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .B1(_3510_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_2275_));
 sky130_fd_sc_hd__nor2_1 _5945_ (.A(_2274_),
    .B(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(_0322_),
    .B(_0639_),
    .Y(_2277_));
 sky130_fd_sc_hd__nand2_1 _5947_ (.A(_0327_),
    .B(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .Y(_2278_));
 sky130_fd_sc_hd__nand2_1 _5948_ (.A(_0332_),
    .B(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .Y(_2279_));
 sky130_fd_sc_hd__nand2_1 _5949_ (.A(_0337_),
    .B(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .Y(_2280_));
 sky130_fd_sc_hd__and4_1 _5950_ (.A(_2277_),
    .B(_2278_),
    .C(_2279_),
    .D(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__and4_1 _5951_ (.A(_2271_),
    .B(_2273_),
    .C(_2276_),
    .D(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__and4_1 _5952_ (.A(_2240_),
    .B(_2254_),
    .C(_2267_),
    .D(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__nor2_1 _5953_ (.A(_3488_),
    .B(_0350_),
    .Y(_2284_));
 sky130_fd_sc_hd__a22o_1 _5954_ (.A1(_0353_),
    .A2(_3497_),
    .B1(_0355_),
    .B2(_0701_),
    .X(_2285_));
 sky130_fd_sc_hd__a211oi_1 _5955_ (.A1(_0796_),
    .A2(_0347_),
    .B1(_2284_),
    .C1(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_0369_),
    .B(_3205_),
    .Y(_2287_));
 sky130_fd_sc_hd__o21ai_1 _5957_ (.A1(_0383_),
    .A2(_0366_),
    .B1(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__a221oi_1 _5958_ (.A1(_3208_),
    .A2(_0360_),
    .B1(_0634_),
    .B2(_0363_),
    .C1(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__o22ai_1 _5959_ (.A1(_0855_),
    .A2(_0381_),
    .B1(_1002_),
    .B2(_0384_),
    .Y(_2290_));
 sky130_fd_sc_hd__a221oi_1 _5960_ (.A1(_0324_),
    .A2(_0375_),
    .B1(_0708_),
    .B2(_0378_),
    .C1(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__nand2_1 _5961_ (.A(_0398_),
    .B(_3482_),
    .Y(_2292_));
 sky130_fd_sc_hd__o21ai_1 _5962_ (.A1(_0697_),
    .A2(_0395_),
    .B1(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__a221oi_1 _5963_ (.A1(_0695_),
    .A2(_0389_),
    .B1(_3476_),
    .B2(_0392_),
    .C1(_2293_),
    .Y(_2294_));
 sky130_fd_sc_hd__and4_1 _5964_ (.A(_2286_),
    .B(_2289_),
    .C(_2291_),
    .D(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_0411_),
    .B(_3189_),
    .Y(_2296_));
 sky130_fd_sc_hd__nand2_1 _5966_ (.A(_0416_),
    .B(_3195_),
    .Y(_2297_));
 sky130_fd_sc_hd__or2_1 _5967_ (.A(_1291_),
    .B(_0421_),
    .X(_2298_));
 sky130_fd_sc_hd__o2111a_1 _5968_ (.A1(_0380_),
    .A2(_0408_),
    .B1(_2296_),
    .C1(_2297_),
    .D1(_2298_),
    .X(_2299_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(_0429_),
    .B(_3163_),
    .Y(_2300_));
 sky130_fd_sc_hd__nand2_1 _5970_ (.A(_0433_),
    .B(_3171_),
    .Y(_2301_));
 sky130_fd_sc_hd__or2_1 _5971_ (.A(_0877_),
    .B(_0438_),
    .X(_2302_));
 sky130_fd_sc_hd__o2111a_1 _5972_ (.A1(_1161_),
    .A2(_0426_),
    .B1(_2300_),
    .C1(_2301_),
    .D1(_2302_),
    .X(_2303_));
 sky130_fd_sc_hd__nand2_1 _5973_ (.A(_0450_),
    .B(_3152_),
    .Y(_2304_));
 sky130_fd_sc_hd__nand2_1 _5974_ (.A(_0455_),
    .B(_0733_),
    .Y(_2305_));
 sky130_fd_sc_hd__nand2_1 _5975_ (.A(_2304_),
    .B(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__a221oi_1 _5976_ (.A1(_0731_),
    .A2(_0444_),
    .B1(_0446_),
    .B2(_0418_),
    .C1(_2306_),
    .Y(_2307_));
 sky130_fd_sc_hd__nand2_1 _5977_ (.A(_0470_),
    .B(_3180_),
    .Y(_2308_));
 sky130_fd_sc_hd__nand2_1 _5978_ (.A(_0474_),
    .B(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_2309_));
 sky130_fd_sc_hd__nand2_1 _5979_ (.A(_2308_),
    .B(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__a221oi_1 _5980_ (.A1(_3183_),
    .A2(_0463_),
    .B1(_3186_),
    .B2(_0467_),
    .C1(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__and4_1 _5981_ (.A(_2299_),
    .B(_2303_),
    .C(_2307_),
    .D(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__nand2_1 _5982_ (.A(_2295_),
    .B(_2312_),
    .Y(_2313_));
 sky130_fd_sc_hd__nand2_1 _5983_ (.A(_0488_),
    .B(_0448_),
    .Y(_2314_));
 sky130_fd_sc_hd__o21ai_1 _5984_ (.A1(_1334_),
    .A2(_0485_),
    .B1(_2314_),
    .Y(_2315_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(_0498_),
    .B(_0442_),
    .Y(_2316_));
 sky130_fd_sc_hd__nand2_1 _5986_ (.A(_0502_),
    .B(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_2317_));
 sky130_fd_sc_hd__nand2_1 _5987_ (.A(_2316_),
    .B(_2317_),
    .Y(_2318_));
 sky130_fd_sc_hd__a221oi_1 _5988_ (.A1(_0919_),
    .A2(_0493_),
    .B1(_0495_),
    .B2(_0534_),
    .C1(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__nand2_1 _5989_ (.A(_0508_),
    .B(_0452_),
    .Y(_2320_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(_0513_),
    .B(_0746_),
    .Y(_2321_));
 sky130_fd_sc_hd__and4b_1 _5991_ (.A_N(_2315_),
    .B(_2319_),
    .C(_2320_),
    .D(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__o22ai_1 _5992_ (.A1(_0437_),
    .A2(_0527_),
    .B1(_0743_),
    .B2(_0530_),
    .Y(_2323_));
 sky130_fd_sc_hd__a221oi_1 _5993_ (.A1(_0741_),
    .A2(_0520_),
    .B1(_0894_),
    .B2(_0524_),
    .C1(_2323_),
    .Y(_2324_));
 sky130_fd_sc_hd__o22ai_1 _5994_ (.A1(_0892_),
    .A2(_0543_),
    .B1(_1037_),
    .B2(_0546_),
    .Y(_2325_));
 sky130_fd_sc_hd__a221oi_1 _5995_ (.A1(_0465_),
    .A2(_0536_),
    .B1(_0413_),
    .B2(_0540_),
    .C1(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__and3_1 _5996_ (.A(_2322_),
    .B(_2324_),
    .C(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__nand2_1 _5997_ (.A(_0562_),
    .B(_1073_),
    .Y(_2328_));
 sky130_fd_sc_hd__nand2_1 _5998_ (.A(_0567_),
    .B(_0932_),
    .Y(_2329_));
 sky130_fd_sc_hd__nand2_1 _5999_ (.A(_2328_),
    .B(_2329_),
    .Y(_2330_));
 sky130_fd_sc_hd__a221oi_1 _6000_ (.A1(_1210_),
    .A2(_0555_),
    .B1(_1055_),
    .B2(_0559_),
    .C1(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__nand2_1 _6001_ (.A(_0582_),
    .B(_0518_),
    .Y(_2332_));
 sky130_fd_sc_hd__nand2_1 _6002_ (.A(_0587_),
    .B(_0916_),
    .Y(_2333_));
 sky130_fd_sc_hd__nand2_1 _6003_ (.A(_2332_),
    .B(_2333_),
    .Y(_2334_));
 sky130_fd_sc_hd__a221oi_1 _6004_ (.A1(_0522_),
    .A2(_0575_),
    .B1(_0768_),
    .B2(_0579_),
    .C1(_2334_),
    .Y(_2335_));
 sky130_fd_sc_hd__nand2_1 _6005_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_2336_));
 sky130_fd_sc_hd__o21ai_1 _6006_ (.A1(_1219_),
    .A2(_0602_),
    .B1(_2336_),
    .Y(_2337_));
 sky130_fd_sc_hd__a221oi_1 _6007_ (.A1(_0577_),
    .A2(_0595_),
    .B1(_0781_),
    .B2(_0599_),
    .C1(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__o22ai_1 _6008_ (.A1(_0481_),
    .A2(_0620_),
    .B1(_0757_),
    .B2(_0623_),
    .Y(_2339_));
 sky130_fd_sc_hd__a221oi_1 _6009_ (.A1(_0515_),
    .A2(_0613_),
    .B1(_0765_),
    .B2(_0617_),
    .C1(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__and4_1 _6010_ (.A(_2331_),
    .B(_2335_),
    .C(_2338_),
    .D(_2340_),
    .X(_2341_));
 sky130_fd_sc_hd__nand2_1 _6011_ (.A(_2327_),
    .B(_2341_),
    .Y(_2342_));
 sky130_fd_sc_hd__nor2_1 _6012_ (.A(_2313_),
    .B(_2342_),
    .Y(_2343_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(_0632_),
    .B(_0865_),
    .Y(_2344_));
 sky130_fd_sc_hd__nand3_1 _6014_ (.A(_2283_),
    .B(_2343_),
    .C(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__nor2_1 _6015_ (.A(_3149_),
    .B(_2345_),
    .Y(_2346_));
 sky130_fd_sc_hd__nor2_1 _6016_ (.A(_2226_),
    .B(_2346_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _6017_ (.A1(_3150_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .B1(_3161_),
    .Y(_2347_));
 sky130_fd_sc_hd__nand2_1 _6018_ (.A(_3236_),
    .B(_0844_),
    .Y(_2348_));
 sky130_fd_sc_hd__nand2_1 _6019_ (.A(_3244_),
    .B(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .Y(_2349_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(_2348_),
    .B(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__a221oi_1 _6021_ (.A1(_0991_),
    .A2(_3222_),
    .B1(_1130_),
    .B2(_3228_),
    .C1(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__nand2_1 _6022_ (.A(_3262_),
    .B(_3453_),
    .Y(_2352_));
 sky130_fd_sc_hd__nand2_1 _6023_ (.A(_3269_),
    .B(_3449_),
    .Y(_2353_));
 sky130_fd_sc_hd__nand2_1 _6024_ (.A(_2352_),
    .B(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__a221oi_1 _6025_ (.A1(_3414_),
    .A2(_3253_),
    .B1(_3418_),
    .B2(_3257_),
    .C1(_2354_),
    .Y(_2355_));
 sky130_fd_sc_hd__nand2_1 _6026_ (.A(_3294_),
    .B(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .Y(_2356_));
 sky130_fd_sc_hd__o21ai_1 _6027_ (.A1(_1499_),
    .A2(_3290_),
    .B1(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__a221oi_1 _6028_ (.A1(_3250_),
    .A2(_3280_),
    .B1(_3285_),
    .B2(_3255_),
    .C1(_2357_),
    .Y(_2358_));
 sky130_fd_sc_hd__o22ai_1 _6029_ (.A1(_0676_),
    .A2(_3313_),
    .B1(_0837_),
    .B2(_3317_),
    .Y(_2359_));
 sky130_fd_sc_hd__a221oi_1 _6030_ (.A1(_0675_),
    .A2(_3304_),
    .B1(_0836_),
    .B2(_3309_),
    .C1(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__and4_1 _6031_ (.A(_2351_),
    .B(_2355_),
    .C(_2358_),
    .D(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__nand2_1 _6032_ (.A(_3334_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_2362_));
 sky130_fd_sc_hd__o21ai_1 _6033_ (.A1(_1219_),
    .A2(_3122_),
    .B1(_2362_),
    .Y(_2363_));
 sky130_fd_sc_hd__a221oi_1 _6034_ (.A1(_0611_),
    .A2(_3325_),
    .B1(_0615_),
    .B2(_3329_),
    .C1(_2363_),
    .Y(_2364_));
 sky130_fd_sc_hd__nand2_1 _6035_ (.A(_3352_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_2365_));
 sky130_fd_sc_hd__o21ai_1 _6036_ (.A1(_1346_),
    .A2(_3349_),
    .B1(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__a221oi_1 _6037_ (.A1(_0593_),
    .A2(_3342_),
    .B1(_0597_),
    .B2(_3346_),
    .C1(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__nand2_1 _6038_ (.A(_3370_),
    .B(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .Y(_2368_));
 sky130_fd_sc_hd__o21ai_1 _6039_ (.A1(_1506_),
    .A2(_3367_),
    .B1(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__a221oi_1 _6040_ (.A1(_0818_),
    .A2(_3360_),
    .B1(_0607_),
    .B2(_3364_),
    .C1(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__nand2_1 _6041_ (.A(_3385_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_2371_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_3389_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_2372_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(_2371_),
    .B(_2372_),
    .Y(_2373_));
 sky130_fd_sc_hd__a221oi_2 _6044_ (.A1(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .A2(_3378_),
    .B1(_0927_),
    .B2(_3382_),
    .C1(_2373_),
    .Y(_2374_));
 sky130_fd_sc_hd__and4_1 _6045_ (.A(_2364_),
    .B(_2367_),
    .C(_2370_),
    .D(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__o22ai_1 _6046_ (.A1(_0827_),
    .A2(_3407_),
    .B1(_0976_),
    .B2(_3410_),
    .Y(_2376_));
 sky130_fd_sc_hd__a221oi_1 _6047_ (.A1(_3340_),
    .A2(_3400_),
    .B1(_3344_),
    .B2(_3404_),
    .C1(_2376_),
    .Y(_2377_));
 sky130_fd_sc_hd__nand2_1 _6048_ (.A(_3426_),
    .B(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .Y(_2378_));
 sky130_fd_sc_hd__o21ai_1 _6049_ (.A1(_1378_),
    .A2(_3423_),
    .B1(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__a221oi_1 _6050_ (.A1(_3376_),
    .A2(_3416_),
    .B1(_3380_),
    .B2(_3420_),
    .C1(_2379_),
    .Y(_2380_));
 sky130_fd_sc_hd__nand2_1 _6051_ (.A(_3444_),
    .B(_3372_),
    .Y(_2381_));
 sky130_fd_sc_hd__o21ai_1 _6052_ (.A1(_3366_),
    .A2(_3441_),
    .B1(_2381_),
    .Y(_2382_));
 sky130_fd_sc_hd__a221oi_1 _6053_ (.A1(_3428_),
    .A2(_3434_),
    .B1(_3437_),
    .B2(_0679_),
    .C1(_2382_),
    .Y(_2383_));
 sky130_fd_sc_hd__nand2_1 _6054_ (.A(_3458_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_2384_));
 sky130_fd_sc_hd__nand2_1 _6055_ (.A(_3462_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_2385_));
 sky130_fd_sc_hd__nand2_1 _6056_ (.A(_2384_),
    .B(_2385_),
    .Y(_2386_));
 sky130_fd_sc_hd__a221oi_1 _6057_ (.A1(_0823_),
    .A2(_3451_),
    .B1(_0972_),
    .B2(_3455_),
    .C1(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__and4_1 _6058_ (.A(_2377_),
    .B(_2380_),
    .C(_2383_),
    .D(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__nand2_1 _6059_ (.A(_3474_),
    .B(_3246_),
    .Y(_2389_));
 sky130_fd_sc_hd__nand2_1 _6060_ (.A(_3479_),
    .B(_0648_),
    .Y(_2390_));
 sky130_fd_sc_hd__or2_1 _6061_ (.A(_0960_),
    .B(_3484_),
    .X(_2391_));
 sky130_fd_sc_hd__o2111a_1 _6062_ (.A1(_0649_),
    .A2(_3471_),
    .B1(_2389_),
    .C1(_2390_),
    .D1(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__nand2_1 _6063_ (.A(_3495_),
    .B(_3287_),
    .Y(_2393_));
 sky130_fd_sc_hd__o221a_1 _6064_ (.A1(_1007_),
    .A2(_3489_),
    .B1(_0861_),
    .B2(_3492_),
    .C1(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__o22ai_1 _6065_ (.A1(_0653_),
    .A2(_3501_),
    .B1(_0814_),
    .B2(_3504_),
    .Y(_2395_));
 sky130_fd_sc_hd__a22o_1 _6066_ (.A1(_3507_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .B1(_3510_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_2396_));
 sky130_fd_sc_hd__nor2_1 _6067_ (.A(_2395_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__nand2_1 _6068_ (.A(_0322_),
    .B(_0801_),
    .Y(_2398_));
 sky130_fd_sc_hd__nand2_1 _6069_ (.A(_0327_),
    .B(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .Y(_2399_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_0332_),
    .B(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .Y(_2400_));
 sky130_fd_sc_hd__nand2_1 _6071_ (.A(_0337_),
    .B(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .Y(_2401_));
 sky130_fd_sc_hd__and4_1 _6072_ (.A(_2398_),
    .B(_2399_),
    .C(_2400_),
    .D(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__and4_1 _6073_ (.A(_2392_),
    .B(_2394_),
    .C(_2397_),
    .D(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__and4_1 _6074_ (.A(_2361_),
    .B(_2375_),
    .C(_2388_),
    .D(_2403_),
    .X(_2404_));
 sky130_fd_sc_hd__nor2_1 _6075_ (.A(_0700_),
    .B(_0350_),
    .Y(_2405_));
 sky130_fd_sc_hd__a22o_1 _6076_ (.A1(_0353_),
    .A2(_0701_),
    .B1(_0355_),
    .B2(_0695_),
    .X(_2406_));
 sky130_fd_sc_hd__a211oi_1 _6077_ (.A1(_0947_),
    .A2(_0347_),
    .B1(_2405_),
    .C1(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__nand2_1 _6078_ (.A(_0369_),
    .B(_3208_),
    .Y(_2408_));
 sky130_fd_sc_hd__o21ai_1 _6079_ (.A1(_0724_),
    .A2(_0366_),
    .B1(_2408_),
    .Y(_2409_));
 sky130_fd_sc_hd__a221oi_1 _6080_ (.A1(_0634_),
    .A2(_0360_),
    .B1(_0796_),
    .B2(_0363_),
    .C1(_2409_),
    .Y(_2410_));
 sky130_fd_sc_hd__o22ai_1 _6081_ (.A1(_1002_),
    .A2(_0381_),
    .B1(_1141_),
    .B2(_0384_),
    .Y(_2411_));
 sky130_fd_sc_hd__a221oi_1 _6082_ (.A1(_0708_),
    .A2(_0375_),
    .B1(_0865_),
    .B2(_0378_),
    .C1(_2411_),
    .Y(_2412_));
 sky130_fd_sc_hd__nand2_1 _6083_ (.A(_0398_),
    .B(_0339_),
    .Y(_2413_));
 sky130_fd_sc_hd__o21ai_1 _6084_ (.A1(_0855_),
    .A2(_0395_),
    .B1(_2413_),
    .Y(_2414_));
 sky130_fd_sc_hd__a221oi_1 _6085_ (.A1(_3476_),
    .A2(_0389_),
    .B1(_3482_),
    .B2(_0392_),
    .C1(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__and4_1 _6086_ (.A(_2407_),
    .B(_2410_),
    .C(_2412_),
    .D(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__nand2_1 _6087_ (.A(_0411_),
    .B(_3192_),
    .Y(_2417_));
 sky130_fd_sc_hd__nand2_1 _6088_ (.A(_0416_),
    .B(_3199_),
    .Y(_2418_));
 sky130_fd_sc_hd__or2_1 _6089_ (.A(_0394_),
    .B(_0421_),
    .X(_2419_));
 sky130_fd_sc_hd__o2111a_1 _6090_ (.A1(_0383_),
    .A2(_0408_),
    .B1(_2417_),
    .C1(_2418_),
    .D1(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__nand2_1 _6091_ (.A(_0429_),
    .B(_3168_),
    .Y(_2421_));
 sky130_fd_sc_hd__nand2_1 _6092_ (.A(_0433_),
    .B(_3174_),
    .Y(_2422_));
 sky130_fd_sc_hd__or2_1 _6093_ (.A(_1022_),
    .B(_0438_),
    .X(_2423_));
 sky130_fd_sc_hd__o2111a_1 _6094_ (.A1(_0349_),
    .A2(_0426_),
    .B1(_2421_),
    .C1(_2422_),
    .D1(_2423_),
    .X(_2424_));
 sky130_fd_sc_hd__nand2_1 _6095_ (.A(_0450_),
    .B(_3163_),
    .Y(_2425_));
 sky130_fd_sc_hd__nand2_1 _6096_ (.A(_0455_),
    .B(_3152_),
    .Y(_2426_));
 sky130_fd_sc_hd__nand2_1 _6097_ (.A(_2425_),
    .B(_2426_),
    .Y(_2427_));
 sky130_fd_sc_hd__a221oi_1 _6098_ (.A1(_0418_),
    .A2(_0444_),
    .B1(_0446_),
    .B2(_0733_),
    .C1(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__nand2_1 _6099_ (.A(_0470_),
    .B(_3183_),
    .Y(_2429_));
 sky130_fd_sc_hd__nand2_1 _6100_ (.A(_0474_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_2430_));
 sky130_fd_sc_hd__nand2_1 _6101_ (.A(_2429_),
    .B(_2430_),
    .Y(_2431_));
 sky130_fd_sc_hd__a221oi_1 _6102_ (.A1(_3186_),
    .A2(_0463_),
    .B1(_3189_),
    .B2(_0467_),
    .C1(_2431_),
    .Y(_2432_));
 sky130_fd_sc_hd__and4_1 _6103_ (.A(_2420_),
    .B(_2424_),
    .C(_2428_),
    .D(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__nand2_1 _6104_ (.A(_2416_),
    .B(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__nand2_1 _6105_ (.A(_0488_),
    .B(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .Y(_2435_));
 sky130_fd_sc_hd__o21ai_1 _6106_ (.A1(_1462_),
    .A2(_0485_),
    .B1(_2435_),
    .Y(_2436_));
 sky130_fd_sc_hd__nand2_1 _6107_ (.A(_0498_),
    .B(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_2437_));
 sky130_fd_sc_hd__nand2_1 _6108_ (.A(_0502_),
    .B(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_2438_));
 sky130_fd_sc_hd__nand2_1 _6109_ (.A(_2437_),
    .B(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__a221oi_1 _6110_ (.A1(_0534_),
    .A2(_0493_),
    .B1(_0495_),
    .B2(_0538_),
    .C1(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_0508_),
    .B(_0746_),
    .Y(_2441_));
 sky130_fd_sc_hd__nand2_1 _6112_ (.A(_0513_),
    .B(_0739_),
    .Y(_2442_));
 sky130_fd_sc_hd__and4b_1 _6113_ (.A_N(_2436_),
    .B(_2440_),
    .C(_2441_),
    .D(_2442_),
    .X(_2443_));
 sky130_fd_sc_hd__o22ai_1 _6114_ (.A1(_0743_),
    .A2(_0527_),
    .B1(_0425_),
    .B2(_0530_),
    .Y(_2444_));
 sky130_fd_sc_hd__a221oi_1 _6115_ (.A1(_0894_),
    .A2(_0520_),
    .B1(_1039_),
    .B2(_0524_),
    .C1(_2444_),
    .Y(_2445_));
 sky130_fd_sc_hd__o22ai_1 _6116_ (.A1(_1037_),
    .A2(_0543_),
    .B1(_1175_),
    .B2(_0546_),
    .Y(_2446_));
 sky130_fd_sc_hd__a221oi_1 _6117_ (.A1(_0413_),
    .A2(_0536_),
    .B1(_0731_),
    .B2(_0540_),
    .C1(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__and3_1 _6118_ (.A(_2443_),
    .B(_2445_),
    .C(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__nand2_1 _6119_ (.A(_0562_),
    .B(_1210_),
    .Y(_2449_));
 sky130_fd_sc_hd__nand2_1 _6120_ (.A(_0567_),
    .B(_1073_),
    .Y(_2450_));
 sky130_fd_sc_hd__nand2_1 _6121_ (.A(_2449_),
    .B(_2450_),
    .Y(_2451_));
 sky130_fd_sc_hd__a221oi_1 _6122_ (.A1(_1055_),
    .A2(_0555_),
    .B1(_1192_),
    .B2(_0559_),
    .C1(_2451_),
    .Y(_2452_));
 sky130_fd_sc_hd__nand2_1 _6123_ (.A(_0582_),
    .B(_0522_),
    .Y(_2453_));
 sky130_fd_sc_hd__nand2_1 _6124_ (.A(_0587_),
    .B(_0518_),
    .Y(_2454_));
 sky130_fd_sc_hd__nand2_1 _6125_ (.A(_2453_),
    .B(_2454_),
    .Y(_2455_));
 sky130_fd_sc_hd__a221oi_1 _6126_ (.A1(_0768_),
    .A2(_0575_),
    .B1(_0919_),
    .B2(_0579_),
    .C1(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hd__nand2_1 _6127_ (.A(_0605_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_2457_));
 sky130_fd_sc_hd__o21ai_1 _6128_ (.A1(_1350_),
    .A2(_0602_),
    .B1(_2457_),
    .Y(_2458_));
 sky130_fd_sc_hd__a221oi_1 _6129_ (.A1(_0781_),
    .A2(_0595_),
    .B1(_0932_),
    .B2(_0599_),
    .C1(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__o22ai_1 _6130_ (.A1(_0757_),
    .A2(_0620_),
    .B1(_0908_),
    .B2(_0623_),
    .Y(_2460_));
 sky130_fd_sc_hd__a221oi_1 _6131_ (.A1(_0765_),
    .A2(_0613_),
    .B1(_0916_),
    .B2(_0617_),
    .C1(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__and4_1 _6132_ (.A(_2452_),
    .B(_2456_),
    .C(_2459_),
    .D(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__nand2_1 _6133_ (.A(_2448_),
    .B(_2462_),
    .Y(_2463_));
 sky130_fd_sc_hd__nor2_1 _6134_ (.A(_2434_),
    .B(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__nand2_1 _6135_ (.A(_0632_),
    .B(_3509_),
    .Y(_2465_));
 sky130_fd_sc_hd__nand3_1 _6136_ (.A(_2404_),
    .B(_2464_),
    .C(_2465_),
    .Y(_2466_));
 sky130_fd_sc_hd__nor2_1 _6137_ (.A(_3149_),
    .B(_2466_),
    .Y(_2467_));
 sky130_fd_sc_hd__nor2_1 _6138_ (.A(_2347_),
    .B(_2467_),
    .Y(_0283_));
 sky130_fd_sc_hd__or4b_1 _6139_ (.A(net47),
    .B(_3124_),
    .C(_3125_),
    .D_N(_3156_),
    .X(_2468_));
 sky130_fd_sc_hd__buf_2 _6140_ (.A(_2468_),
    .X(_2469_));
 sky130_fd_sc_hd__clkbuf_4 _6141_ (.A(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__buf_4 _6142_ (.A(_3156_),
    .X(_2471_));
 sky130_fd_sc_hd__a31o_1 _6143_ (.A1(_2471_),
    .A2(\egd_top.BitStream_buffer.buffer_index[5] ),
    .A3(\egd_top.BitStream_buffer.buffer_index[4] ),
    .B1(_3132_),
    .X(_2472_));
 sky130_fd_sc_hd__a21oi_1 _6144_ (.A1(_2470_),
    .A2(_2472_),
    .B1(_3090_),
    .Y(_0282_));
 sky130_fd_sc_hd__or2_1 _6145_ (.A(_3124_),
    .B(_2471_),
    .X(_2473_));
 sky130_fd_sc_hd__nor2_2 _6146_ (.A(net44),
    .B(net46),
    .Y(_2474_));
 sky130_fd_sc_hd__nor2_2 _6147_ (.A(net45),
    .B(_3124_),
    .Y(_2475_));
 sky130_fd_sc_hd__o21ai_1 _6148_ (.A1(_2474_),
    .A2(_2475_),
    .B1(_2471_),
    .Y(_2476_));
 sky130_fd_sc_hd__a21oi_1 _6149_ (.A1(_2473_),
    .A2(_2476_),
    .B1(_3089_),
    .Y(_0281_));
 sky130_fd_sc_hd__or2_1 _6150_ (.A(_3125_),
    .B(_2471_),
    .X(_2477_));
 sky130_fd_sc_hd__nand2_1 _6151_ (.A(_2471_),
    .B(_3125_),
    .Y(_2478_));
 sky130_fd_sc_hd__a21oi_1 _6152_ (.A1(_2477_),
    .A2(_2478_),
    .B1(_3089_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_4 _6153_ (.A(_2471_),
    .B(_3133_),
    .Y(_2479_));
 sky130_fd_sc_hd__clkbuf_4 _6154_ (.A(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__mux2_1 _6155_ (.A0(net7),
    .A1(_0634_),
    .S(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__and2_1 _6156_ (.A(_2481_),
    .B(_3197_),
    .X(_2482_));
 sky130_fd_sc_hd__clkbuf_1 _6157_ (.A(_2482_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _6158_ (.A0(net6),
    .A1(_0796_),
    .S(_2480_),
    .X(_2483_));
 sky130_fd_sc_hd__and2_1 _6159_ (.A(_2483_),
    .B(_3197_),
    .X(_2484_));
 sky130_fd_sc_hd__clkbuf_1 _6160_ (.A(_2484_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _6161_ (.A0(net5),
    .A1(_0947_),
    .S(_2480_),
    .X(_2485_));
 sky130_fd_sc_hd__and2_1 _6162_ (.A(_2485_),
    .B(_3197_),
    .X(_2486_));
 sky130_fd_sc_hd__clkbuf_1 _6163_ (.A(_2486_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _6164_ (.A0(net4),
    .A1(_3497_),
    .S(_2480_),
    .X(_2487_));
 sky130_fd_sc_hd__and2_1 _6165_ (.A(_2487_),
    .B(_3197_),
    .X(_2488_));
 sky130_fd_sc_hd__clkbuf_1 _6166_ (.A(_2488_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _6167_ (.A0(net3),
    .A1(_0701_),
    .S(_2480_),
    .X(_2489_));
 sky130_fd_sc_hd__and2_1 _6168_ (.A(_2489_),
    .B(_3197_),
    .X(_2490_));
 sky130_fd_sc_hd__clkbuf_1 _6169_ (.A(_2490_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _6170_ (.A0(net2),
    .A1(_0695_),
    .S(_2480_),
    .X(_2491_));
 sky130_fd_sc_hd__buf_8 _6171_ (.A(_3165_),
    .X(_2492_));
 sky130_fd_sc_hd__and2_1 _6172_ (.A(_2491_),
    .B(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__clkbuf_1 _6173_ (.A(_2493_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _6174_ (.A0(net16),
    .A1(_3476_),
    .S(_2480_),
    .X(_2494_));
 sky130_fd_sc_hd__and2_1 _6175_ (.A(_2492_),
    .B(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__clkbuf_1 _6176_ (.A(_2495_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _6177_ (.A0(net15),
    .A1(_3482_),
    .S(_2480_),
    .X(_2496_));
 sky130_fd_sc_hd__and2_4 _6178_ (.A(_2496_),
    .B(_2492_),
    .X(_2497_));
 sky130_fd_sc_hd__clkbuf_1 _6179_ (.A(_2497_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _6180_ (.A0(net14),
    .A1(_0339_),
    .S(_2480_),
    .X(_2498_));
 sky130_fd_sc_hd__and2_4 _6181_ (.A(_2498_),
    .B(_2492_),
    .X(_2499_));
 sky130_fd_sc_hd__clkbuf_1 _6182_ (.A(_2499_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _6183_ (.A0(net13),
    .A1(_0329_),
    .S(_2480_),
    .X(_2500_));
 sky130_fd_sc_hd__and2_1 _6184_ (.A(_2492_),
    .B(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__clkbuf_1 _6185_ (.A(_2501_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _6186_ (.A0(net12),
    .A1(_0334_),
    .S(_2479_),
    .X(_2502_));
 sky130_fd_sc_hd__and2_1 _6187_ (.A(_2502_),
    .B(_2492_),
    .X(_2503_));
 sky130_fd_sc_hd__clkbuf_1 _6188_ (.A(_2503_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _6189_ (.A0(net11),
    .A1(_0324_),
    .S(_2479_),
    .X(_2504_));
 sky130_fd_sc_hd__and2_1 _6190_ (.A(_2492_),
    .B(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__clkbuf_1 _6191_ (.A(_2505_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _6192_ (.A0(net10),
    .A1(_0708_),
    .S(_2479_),
    .X(_2506_));
 sky130_fd_sc_hd__and2_4 _6193_ (.A(_2506_),
    .B(_2492_),
    .X(_2507_));
 sky130_fd_sc_hd__clkbuf_1 _6194_ (.A(_2507_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _6195_ (.A0(net9),
    .A1(_0865_),
    .S(_2479_),
    .X(_2508_));
 sky130_fd_sc_hd__and2_1 _6196_ (.A(_2492_),
    .B(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__clkbuf_1 _6197_ (.A(_2509_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _6198_ (.A0(net8),
    .A1(_3509_),
    .S(_2479_),
    .X(_2510_));
 sky130_fd_sc_hd__and2_1 _6199_ (.A(_2492_),
    .B(_2510_),
    .X(_2511_));
 sky130_fd_sc_hd__clkbuf_1 _6200_ (.A(_2511_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _6201_ (.A0(net1),
    .A1(_3512_),
    .S(_2479_),
    .X(_2512_));
 sky130_fd_sc_hd__buf_8 _6202_ (.A(_3165_),
    .X(_2513_));
 sky130_fd_sc_hd__and2_1 _6203_ (.A(_2512_),
    .B(_2513_),
    .X(_2514_));
 sky130_fd_sc_hd__clkbuf_1 _6204_ (.A(_2514_),
    .X(_0264_));
 sky130_fd_sc_hd__nand3_4 _6205_ (.A(_2471_),
    .B(_3132_),
    .C(_2474_),
    .Y(_2515_));
 sky130_fd_sc_hd__clkbuf_4 _6206_ (.A(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__mux2_1 _6207_ (.A0(net7),
    .A1(_3275_),
    .S(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__and2_1 _6208_ (.A(_2517_),
    .B(_2513_),
    .X(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _6209_ (.A(_2518_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _6210_ (.A0(net6),
    .A1(_3287_),
    .S(_2516_),
    .X(_2519_));
 sky130_fd_sc_hd__and2_1 _6211_ (.A(_2519_),
    .B(_2513_),
    .X(_2520_));
 sky130_fd_sc_hd__clkbuf_1 _6212_ (.A(_2520_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _6213_ (.A0(net5),
    .A1(_0648_),
    .S(_2516_),
    .X(_2521_));
 sky130_fd_sc_hd__and2_1 _6214_ (.A(_2521_),
    .B(_2513_),
    .X(_2522_));
 sky130_fd_sc_hd__clkbuf_1 _6215_ (.A(_2522_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _6216_ (.A0(net4),
    .A1(_3296_),
    .S(_2516_),
    .X(_2523_));
 sky130_fd_sc_hd__and2_1 _6217_ (.A(_2513_),
    .B(_2523_),
    .X(_2524_));
 sky130_fd_sc_hd__clkbuf_1 _6218_ (.A(_2524_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _6219_ (.A0(net3),
    .A1(_3246_),
    .S(_2516_),
    .X(_2525_));
 sky130_fd_sc_hd__and2_1 _6220_ (.A(_2525_),
    .B(_2513_),
    .X(_2526_));
 sky130_fd_sc_hd__clkbuf_1 _6221_ (.A(_2526_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _6222_ (.A0(net2),
    .A1(_3238_),
    .S(_2516_),
    .X(_2527_));
 sky130_fd_sc_hd__and2_1 _6223_ (.A(_2513_),
    .B(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__clkbuf_1 _6224_ (.A(_2528_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _6225_ (.A0(net16),
    .A1(_3213_),
    .S(_2516_),
    .X(_2529_));
 sky130_fd_sc_hd__and2_1 _6226_ (.A(_2513_),
    .B(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__clkbuf_1 _6227_ (.A(_2530_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _6228_ (.A0(net15),
    .A1(_3224_),
    .S(_2516_),
    .X(_2531_));
 sky130_fd_sc_hd__and2_1 _6229_ (.A(_2513_),
    .B(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__clkbuf_1 _6230_ (.A(_2532_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _6231_ (.A0(net14),
    .A1(_0639_),
    .S(_2516_),
    .X(_2533_));
 sky130_fd_sc_hd__and2_1 _6232_ (.A(_2513_),
    .B(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__clkbuf_1 _6233_ (.A(_2534_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _6234_ (.A0(net13),
    .A1(_0801_),
    .S(_2516_),
    .X(_2535_));
 sky130_fd_sc_hd__buf_6 _6235_ (.A(_3165_),
    .X(_2536_));
 sky130_fd_sc_hd__and2_1 _6236_ (.A(_2535_),
    .B(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__clkbuf_1 _6237_ (.A(_2537_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _6238_ (.A0(net12),
    .A1(_3300_),
    .S(_2515_),
    .X(_2538_));
 sky130_fd_sc_hd__and2_1 _6239_ (.A(_2538_),
    .B(_2536_),
    .X(_2539_));
 sky130_fd_sc_hd__clkbuf_1 _6240_ (.A(_2539_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _6241_ (.A0(net11),
    .A1(_3306_),
    .S(_2515_),
    .X(_2540_));
 sky130_fd_sc_hd__and2_1 _6242_ (.A(_2540_),
    .B(_2536_),
    .X(_2541_));
 sky130_fd_sc_hd__clkbuf_1 _6243_ (.A(_2541_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _6244_ (.A0(net10),
    .A1(_3271_),
    .S(_2515_),
    .X(_2542_));
 sky130_fd_sc_hd__and2_1 _6245_ (.A(_2542_),
    .B(_2536_),
    .X(_2543_));
 sky130_fd_sc_hd__clkbuf_1 _6246_ (.A(_2543_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _6247_ (.A0(net9),
    .A1(_3264_),
    .S(_2515_),
    .X(_2544_));
 sky130_fd_sc_hd__and2_1 _6248_ (.A(_2544_),
    .B(_2536_),
    .X(_2545_));
 sky130_fd_sc_hd__clkbuf_1 _6249_ (.A(_2545_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _6250_ (.A0(net8),
    .A1(_3250_),
    .S(_2515_),
    .X(_2546_));
 sky130_fd_sc_hd__and2_1 _6251_ (.A(_2546_),
    .B(_2536_),
    .X(_2547_));
 sky130_fd_sc_hd__clkbuf_1 _6252_ (.A(_2547_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _6253_ (.A0(net1),
    .A1(_3255_),
    .S(_2515_),
    .X(_2548_));
 sky130_fd_sc_hd__and2_1 _6254_ (.A(_2548_),
    .B(_2536_),
    .X(_2549_));
 sky130_fd_sc_hd__clkbuf_1 _6255_ (.A(_2549_),
    .X(_0248_));
 sky130_fd_sc_hd__nand3_4 _6256_ (.A(_2471_),
    .B(_3132_),
    .C(_2475_),
    .Y(_2550_));
 sky130_fd_sc_hd__clkbuf_4 _6257_ (.A(_2550_),
    .X(_2551_));
 sky130_fd_sc_hd__mux2_1 _6258_ (.A0(net7),
    .A1(_3432_),
    .S(_2551_),
    .X(_2552_));
 sky130_fd_sc_hd__and2_1 _6259_ (.A(_2552_),
    .B(_2536_),
    .X(_2553_));
 sky130_fd_sc_hd__clkbuf_1 _6260_ (.A(_2553_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _6261_ (.A0(net6),
    .A1(_3439_),
    .S(_2551_),
    .X(_2554_));
 sky130_fd_sc_hd__and2_1 _6262_ (.A(_2554_),
    .B(_2536_),
    .X(_2555_));
 sky130_fd_sc_hd__clkbuf_1 _6263_ (.A(_2555_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _6264_ (.A0(net5),
    .A1(_0683_),
    .S(_2551_),
    .X(_2556_));
 sky130_fd_sc_hd__and2_1 _6265_ (.A(_2556_),
    .B(_2536_),
    .X(_2557_));
 sky130_fd_sc_hd__clkbuf_1 _6266_ (.A(_2557_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _6267_ (.A0(net4),
    .A1(_0844_),
    .S(_2551_),
    .X(_2558_));
 sky130_fd_sc_hd__clkbuf_2 _6268_ (.A(net39),
    .X(_2559_));
 sky130_fd_sc_hd__and2_1 _6269_ (.A(_2558_),
    .B(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__clkbuf_1 _6270_ (.A(_2560_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _6271_ (.A0(net3),
    .A1(_0991_),
    .S(_2551_),
    .X(_2561_));
 sky130_fd_sc_hd__and2_1 _6272_ (.A(_2561_),
    .B(_2559_),
    .X(_2562_));
 sky130_fd_sc_hd__clkbuf_1 _6273_ (.A(_2562_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _6274_ (.A0(net2),
    .A1(_1130_),
    .S(_2551_),
    .X(_2563_));
 sky130_fd_sc_hd__and2_1 _6275_ (.A(_2563_),
    .B(_2559_),
    .X(_2564_));
 sky130_fd_sc_hd__clkbuf_1 _6276_ (.A(_2564_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _6277_ (.A0(net16),
    .A1(_3395_),
    .S(_2551_),
    .X(_2565_));
 sky130_fd_sc_hd__and2_1 _6278_ (.A(_2565_),
    .B(_2559_),
    .X(_2566_));
 sky130_fd_sc_hd__clkbuf_1 _6279_ (.A(_2566_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _6280_ (.A0(net15),
    .A1(_3402_),
    .S(_2551_),
    .X(_2567_));
 sky130_fd_sc_hd__and2_1 _6281_ (.A(_2567_),
    .B(_2559_),
    .X(_2568_));
 sky130_fd_sc_hd__clkbuf_1 _6282_ (.A(_2568_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _6283_ (.A0(net14),
    .A1(_0675_),
    .S(_2551_),
    .X(_2569_));
 sky130_fd_sc_hd__and2_1 _6284_ (.A(_2569_),
    .B(_2559_),
    .X(_2570_));
 sky130_fd_sc_hd__clkbuf_1 _6285_ (.A(_2570_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _6286_ (.A0(net13),
    .A1(_0836_),
    .S(_2551_),
    .X(_2571_));
 sky130_fd_sc_hd__and2_1 _6287_ (.A(_2571_),
    .B(_2559_),
    .X(_2572_));
 sky130_fd_sc_hd__clkbuf_1 _6288_ (.A(_2572_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _6289_ (.A0(net12),
    .A1(_3449_),
    .S(_2550_),
    .X(_2573_));
 sky130_fd_sc_hd__and2_1 _6290_ (.A(_2573_),
    .B(_2559_),
    .X(_2574_));
 sky130_fd_sc_hd__clkbuf_1 _6291_ (.A(_2574_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _6292_ (.A0(net11),
    .A1(_3453_),
    .S(_2550_),
    .X(_2575_));
 sky130_fd_sc_hd__and2_1 _6293_ (.A(_2575_),
    .B(_2559_),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_1 _6294_ (.A(_2576_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _6295_ (.A0(net10),
    .A1(_3414_),
    .S(_2550_),
    .X(_2577_));
 sky130_fd_sc_hd__and2_1 _6296_ (.A(_2577_),
    .B(_2559_),
    .X(_2578_));
 sky130_fd_sc_hd__clkbuf_1 _6297_ (.A(_2578_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _6298_ (.A0(net9),
    .A1(_3418_),
    .S(_2550_),
    .X(_2579_));
 sky130_fd_sc_hd__clkbuf_2 _6299_ (.A(net39),
    .X(_2580_));
 sky130_fd_sc_hd__and2_1 _6300_ (.A(_2579_),
    .B(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__clkbuf_1 _6301_ (.A(_2581_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _6302_ (.A0(net8),
    .A1(_3428_),
    .S(_2550_),
    .X(_2582_));
 sky130_fd_sc_hd__and2_1 _6303_ (.A(_2582_),
    .B(_2580_),
    .X(_2583_));
 sky130_fd_sc_hd__clkbuf_1 _6304_ (.A(_2583_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _6305_ (.A0(net1),
    .A1(_0679_),
    .S(_2550_),
    .X(_2584_));
 sky130_fd_sc_hd__and2_1 _6306_ (.A(_2584_),
    .B(_2580_),
    .X(_2585_));
 sky130_fd_sc_hd__clkbuf_1 _6307_ (.A(_2585_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _6308_ (.A0(net7),
    .A1(_0840_),
    .S(_2470_),
    .X(_2586_));
 sky130_fd_sc_hd__and2_1 _6309_ (.A(_2586_),
    .B(_2580_),
    .X(_2587_));
 sky130_fd_sc_hd__clkbuf_1 _6310_ (.A(_2587_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _6311_ (.A0(net6),
    .A1(_3372_),
    .S(_2470_),
    .X(_2588_));
 sky130_fd_sc_hd__and2_1 _6312_ (.A(_2588_),
    .B(_2580_),
    .X(_2589_));
 sky130_fd_sc_hd__clkbuf_1 _6313_ (.A(_2589_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _6314_ (.A0(net5),
    .A1(_3358_),
    .S(_2470_),
    .X(_2590_));
 sky130_fd_sc_hd__and2_1 _6315_ (.A(_2590_),
    .B(_2580_),
    .X(_2591_));
 sky130_fd_sc_hd__clkbuf_1 _6316_ (.A(_2591_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _6317_ (.A0(net4),
    .A1(_3362_),
    .S(_2470_),
    .X(_2592_));
 sky130_fd_sc_hd__and2_1 _6318_ (.A(_2592_),
    .B(_2580_),
    .X(_2593_));
 sky130_fd_sc_hd__clkbuf_1 _6319_ (.A(_2593_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _6320_ (.A0(net3),
    .A1(_3340_),
    .S(_2470_),
    .X(_2594_));
 sky130_fd_sc_hd__and2_1 _6321_ (.A(_2594_),
    .B(_2580_),
    .X(_2595_));
 sky130_fd_sc_hd__clkbuf_1 _6322_ (.A(_2595_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _6323_ (.A0(net2),
    .A1(_3344_),
    .S(_2470_),
    .X(_2596_));
 sky130_fd_sc_hd__and2_1 _6324_ (.A(_2596_),
    .B(_2580_),
    .X(_2597_));
 sky130_fd_sc_hd__clkbuf_1 _6325_ (.A(_2597_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _6326_ (.A0(net16),
    .A1(_3354_),
    .S(_2470_),
    .X(_2598_));
 sky130_fd_sc_hd__and2_1 _6327_ (.A(_2598_),
    .B(_2580_),
    .X(_2599_));
 sky130_fd_sc_hd__clkbuf_1 _6328_ (.A(_2599_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _6329_ (.A0(net15),
    .A1(_0662_),
    .S(_2470_),
    .X(_2600_));
 sky130_fd_sc_hd__clkbuf_2 _6330_ (.A(net39),
    .X(_2601_));
 sky130_fd_sc_hd__and2_1 _6331_ (.A(_2600_),
    .B(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__clkbuf_1 _6332_ (.A(_2602_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _6333_ (.A0(net14),
    .A1(_0823_),
    .S(_2470_),
    .X(_2603_));
 sky130_fd_sc_hd__and2_1 _6334_ (.A(_2603_),
    .B(_2601_),
    .X(_2604_));
 sky130_fd_sc_hd__clkbuf_1 _6335_ (.A(_2604_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _6336_ (.A0(net13),
    .A1(_0972_),
    .S(_2469_),
    .X(_2605_));
 sky130_fd_sc_hd__and2_1 _6337_ (.A(_2605_),
    .B(_2601_),
    .X(_2606_));
 sky130_fd_sc_hd__clkbuf_1 _6338_ (.A(_2606_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _6339_ (.A0(net12),
    .A1(_3376_),
    .S(_2469_),
    .X(_2607_));
 sky130_fd_sc_hd__and2_1 _6340_ (.A(_2607_),
    .B(_2601_),
    .X(_2608_));
 sky130_fd_sc_hd__clkbuf_1 _6341_ (.A(_2608_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _6342_ (.A0(net11),
    .A1(_3380_),
    .S(_2469_),
    .X(_2609_));
 sky130_fd_sc_hd__and2_1 _6343_ (.A(_2609_),
    .B(_2601_),
    .X(_2610_));
 sky130_fd_sc_hd__clkbuf_1 _6344_ (.A(_2610_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _6345_ (.A0(net10),
    .A1(_3322_),
    .S(_2469_),
    .X(_2611_));
 sky130_fd_sc_hd__and2_1 _6346_ (.A(_2611_),
    .B(_2601_),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_1 _6347_ (.A(_2612_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _6348_ (.A0(net9),
    .A1(_3327_),
    .S(_2469_),
    .X(_2613_));
 sky130_fd_sc_hd__and2_1 _6349_ (.A(_2613_),
    .B(_2601_),
    .X(_2614_));
 sky130_fd_sc_hd__clkbuf_1 _6350_ (.A(_2614_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _6351_ (.A0(net8),
    .A1(_3336_),
    .S(_2469_),
    .X(_2615_));
 sky130_fd_sc_hd__and2_1 _6352_ (.A(_2615_),
    .B(_2601_),
    .X(_2616_));
 sky130_fd_sc_hd__clkbuf_1 _6353_ (.A(_2616_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _6354_ (.A0(net1),
    .A1(_0657_),
    .S(_2469_),
    .X(_2617_));
 sky130_fd_sc_hd__and2_1 _6355_ (.A(_2617_),
    .B(_2601_),
    .X(_2618_));
 sky130_fd_sc_hd__clkbuf_1 _6356_ (.A(_2618_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_4 _6357_ (.A(_2471_),
    .B(_3126_),
    .Y(_2619_));
 sky130_fd_sc_hd__clkbuf_4 _6358_ (.A(_2619_),
    .X(_2620_));
 sky130_fd_sc_hd__mux2_1 _6359_ (.A0(net7),
    .A1(_0818_),
    .S(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__and2_1 _6360_ (.A(_2621_),
    .B(_2601_),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_1 _6361_ (.A(_2622_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _6362_ (.A0(net6),
    .A1(_0607_),
    .S(_2620_),
    .X(_2623_));
 sky130_fd_sc_hd__clkbuf_2 _6363_ (.A(net39),
    .X(_2624_));
 sky130_fd_sc_hd__and2_1 _6364_ (.A(_2623_),
    .B(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__clkbuf_1 _6365_ (.A(_2625_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _6366_ (.A0(net5),
    .A1(_0593_),
    .S(_2620_),
    .X(_2626_));
 sky130_fd_sc_hd__and2_1 _6367_ (.A(_2626_),
    .B(_2624_),
    .X(_2627_));
 sky130_fd_sc_hd__clkbuf_1 _6368_ (.A(_2627_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _6369_ (.A0(net4),
    .A1(_0597_),
    .S(_2620_),
    .X(_2628_));
 sky130_fd_sc_hd__and2_1 _6370_ (.A(_2628_),
    .B(_2624_),
    .X(_2629_));
 sky130_fd_sc_hd__clkbuf_1 _6371_ (.A(_2629_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _6372_ (.A0(net3),
    .A1(_0569_),
    .S(_2620_),
    .X(_2630_));
 sky130_fd_sc_hd__and2_1 _6373_ (.A(_2630_),
    .B(_2624_),
    .X(_2631_));
 sky130_fd_sc_hd__clkbuf_1 _6374_ (.A(_2631_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _6375_ (.A0(net2),
    .A1(_0564_),
    .S(_2620_),
    .X(_2632_));
 sky130_fd_sc_hd__and2_1 _6376_ (.A(_2632_),
    .B(_2624_),
    .X(_2633_));
 sky130_fd_sc_hd__clkbuf_1 _6377_ (.A(_2633_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _6378_ (.A0(net16),
    .A1(_0551_),
    .S(_2620_),
    .X(_2634_));
 sky130_fd_sc_hd__and2_1 _6379_ (.A(_2634_),
    .B(_2624_),
    .X(_2635_));
 sky130_fd_sc_hd__clkbuf_1 _6380_ (.A(_2635_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _6381_ (.A0(net15),
    .A1(_0557_),
    .S(_2620_),
    .X(_2636_));
 sky130_fd_sc_hd__and2_1 _6382_ (.A(_2636_),
    .B(_2624_),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_1 _6383_ (.A(_2637_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _6384_ (.A0(net14),
    .A1(_0776_),
    .S(_2620_),
    .X(_2638_));
 sky130_fd_sc_hd__and2_1 _6385_ (.A(_2638_),
    .B(_2624_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _6386_ (.A(_2639_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _6387_ (.A0(net13),
    .A1(_0927_),
    .S(_2620_),
    .X(_2640_));
 sky130_fd_sc_hd__and2_1 _6388_ (.A(_2640_),
    .B(_2624_),
    .X(_2641_));
 sky130_fd_sc_hd__clkbuf_1 _6389_ (.A(_2641_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _6390_ (.A0(net12),
    .A1(_0611_),
    .S(_2619_),
    .X(_2642_));
 sky130_fd_sc_hd__and2_1 _6391_ (.A(_2642_),
    .B(_2624_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _6392_ (.A(_2643_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _6393_ (.A0(net11),
    .A1(_0615_),
    .S(_2619_),
    .X(_2644_));
 sky130_fd_sc_hd__buf_2 _6394_ (.A(net39),
    .X(_2645_));
 sky130_fd_sc_hd__and2_1 _6395_ (.A(_2644_),
    .B(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__clkbuf_1 _6396_ (.A(_2646_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _6397_ (.A0(net10),
    .A1(_0589_),
    .S(_2619_),
    .X(_2647_));
 sky130_fd_sc_hd__and2_1 _6398_ (.A(_2647_),
    .B(_2645_),
    .X(_2648_));
 sky130_fd_sc_hd__clkbuf_1 _6399_ (.A(_2648_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _6400_ (.A0(net9),
    .A1(_0584_),
    .S(_2619_),
    .X(_2649_));
 sky130_fd_sc_hd__and2_1 _6401_ (.A(_2649_),
    .B(_2645_),
    .X(_2650_));
 sky130_fd_sc_hd__clkbuf_1 _6402_ (.A(_2650_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _6403_ (.A0(net8),
    .A1(_0573_),
    .S(_2619_),
    .X(_2651_));
 sky130_fd_sc_hd__and2_1 _6404_ (.A(_2651_),
    .B(_2645_),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _6405_ (.A(_2652_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _6406_ (.A0(net1),
    .A1(_0577_),
    .S(_2619_),
    .X(_2653_));
 sky130_fd_sc_hd__and2_1 _6407_ (.A(_2653_),
    .B(_2645_),
    .X(_2654_));
 sky130_fd_sc_hd__clkbuf_1 _6408_ (.A(_2654_),
    .X(_0200_));
 sky130_fd_sc_hd__nand3_2 _6409_ (.A(_2471_),
    .B(net42),
    .C(_2475_),
    .Y(_2655_));
 sky130_fd_sc_hd__clkbuf_4 _6410_ (.A(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__mux2_1 _6411_ (.A0(net7),
    .A1(_0442_),
    .S(_2656_),
    .X(_2657_));
 sky130_fd_sc_hd__and2_1 _6412_ (.A(_2657_),
    .B(_2645_),
    .X(_2658_));
 sky130_fd_sc_hd__clkbuf_1 _6413_ (.A(_2658_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _6414_ (.A0(net6),
    .A1(_0448_),
    .S(_2656_),
    .X(_2659_));
 sky130_fd_sc_hd__and2_1 _6415_ (.A(_2659_),
    .B(_2645_),
    .X(_2660_));
 sky130_fd_sc_hd__clkbuf_1 _6416_ (.A(_2660_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _6417_ (.A0(net5),
    .A1(_0457_),
    .S(_2656_),
    .X(_2661_));
 sky130_fd_sc_hd__and2_1 _6418_ (.A(_2661_),
    .B(_2645_),
    .X(_2662_));
 sky130_fd_sc_hd__clkbuf_1 _6419_ (.A(_2662_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _6420_ (.A0(net4),
    .A1(_0452_),
    .S(_2656_),
    .X(_2663_));
 sky130_fd_sc_hd__and2_1 _6421_ (.A(_2663_),
    .B(_2645_),
    .X(_2664_));
 sky130_fd_sc_hd__clkbuf_1 _6422_ (.A(_2664_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _6423_ (.A0(net3),
    .A1(_0746_),
    .S(_2656_),
    .X(_2665_));
 sky130_fd_sc_hd__and2_1 _6424_ (.A(_2665_),
    .B(_2645_),
    .X(_2666_));
 sky130_fd_sc_hd__clkbuf_1 _6425_ (.A(_2666_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _6426_ (.A0(net2),
    .A1(_0739_),
    .S(_2656_),
    .X(_2667_));
 sky130_fd_sc_hd__clkbuf_2 _6427_ (.A(_3079_),
    .X(_2668_));
 sky130_fd_sc_hd__and2_1 _6428_ (.A(_2667_),
    .B(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__clkbuf_1 _6429_ (.A(_2669_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _6430_ (.A0(net16),
    .A1(_0435_),
    .S(_2656_),
    .X(_2670_));
 sky130_fd_sc_hd__and2_1 _6431_ (.A(_2670_),
    .B(_2668_),
    .X(_2671_));
 sky130_fd_sc_hd__clkbuf_1 _6432_ (.A(_2671_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _6433_ (.A0(net15),
    .A1(_0741_),
    .S(_2656_),
    .X(_2672_));
 sky130_fd_sc_hd__and2_1 _6434_ (.A(_2672_),
    .B(_2668_),
    .X(_2673_));
 sky130_fd_sc_hd__clkbuf_1 _6435_ (.A(_2673_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _6436_ (.A0(net14),
    .A1(_0894_),
    .S(_2656_),
    .X(_2674_));
 sky130_fd_sc_hd__and2_1 _6437_ (.A(_2674_),
    .B(_2668_),
    .X(_2675_));
 sky130_fd_sc_hd__clkbuf_1 _6438_ (.A(_2675_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _6439_ (.A0(net13),
    .A1(_1039_),
    .S(_2656_),
    .X(_2676_));
 sky130_fd_sc_hd__and2_1 _6440_ (.A(_2676_),
    .B(_2668_),
    .X(_2677_));
 sky130_fd_sc_hd__clkbuf_1 _6441_ (.A(_2677_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _6442_ (.A0(net12),
    .A1(_0461_),
    .S(net43),
    .X(_2678_));
 sky130_fd_sc_hd__and2_1 _6443_ (.A(_2678_),
    .B(_2668_),
    .X(_2679_));
 sky130_fd_sc_hd__clkbuf_1 _6444_ (.A(_2679_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _6445_ (.A0(net11),
    .A1(_0465_),
    .S(net43),
    .X(_2680_));
 sky130_fd_sc_hd__and2_1 _6446_ (.A(_2680_),
    .B(_2668_),
    .X(_2681_));
 sky130_fd_sc_hd__clkbuf_1 _6447_ (.A(_2681_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _6448_ (.A0(net10),
    .A1(_0413_),
    .S(net43),
    .X(_2682_));
 sky130_fd_sc_hd__and2_1 _6449_ (.A(_2682_),
    .B(_2668_),
    .X(_2683_));
 sky130_fd_sc_hd__clkbuf_1 _6450_ (.A(_2683_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _6451_ (.A0(net9),
    .A1(_0731_),
    .S(net43),
    .X(_2684_));
 sky130_fd_sc_hd__and2_1 _6452_ (.A(_2684_),
    .B(_2668_),
    .X(_2685_));
 sky130_fd_sc_hd__clkbuf_1 _6453_ (.A(_2685_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _6454_ (.A0(net8),
    .A1(_0418_),
    .S(net43),
    .X(_2686_));
 sky130_fd_sc_hd__and2_1 _6455_ (.A(_2686_),
    .B(_2668_),
    .X(_2687_));
 sky130_fd_sc_hd__clkbuf_1 _6456_ (.A(_2687_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _6457_ (.A0(net1),
    .A1(_0733_),
    .S(net43),
    .X(_2688_));
 sky130_fd_sc_hd__buf_2 _6458_ (.A(_3079_),
    .X(_2689_));
 sky130_fd_sc_hd__and2_1 _6459_ (.A(_2688_),
    .B(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__clkbuf_1 _6460_ (.A(_2690_),
    .X(_0184_));
 sky130_fd_sc_hd__nor2_1 _6461_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2691_));
 sky130_fd_sc_hd__nand2_1 _6462_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2692_));
 sky130_fd_sc_hd__o21ai_4 _6463_ (.A1(_2691_),
    .A2(_3113_),
    .B1(_2692_),
    .Y(_2693_));
 sky130_fd_sc_hd__or2_1 _6464_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .X(_2694_));
 sky130_fd_sc_hd__nand2_1 _6465_ (.A(\egd_top.BitStream_buffer.pc_previous[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2695_));
 sky130_fd_sc_hd__a21bo_2 _6466_ (.A1(_2693_),
    .A2(_2694_),
    .B1_N(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__or2_1 _6467_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .X(_2697_));
 sky130_fd_sc_hd__nand2_1 _6468_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2698_));
 sky130_fd_sc_hd__a21bo_2 _6469_ (.A1(_2696_),
    .A2(_2697_),
    .B1_N(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__and3_2 _6470_ (.A(_2699_),
    .B(\egd_top.BitStream_buffer.pc_previous[4] ),
    .C(\egd_top.BitStream_buffer.pc_previous[5] ),
    .X(_2700_));
 sky130_fd_sc_hd__xor2_4 _6471_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .B(_2700_),
    .X(\egd_top.BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nor2_1 _6472_ (.A(_3120_),
    .B(_3090_),
    .Y(_0183_));
 sky130_fd_sc_hd__a21oi_1 _6473_ (.A1(_2699_),
    .A2(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B1(\egd_top.BitStream_buffer.pc_previous[5] ),
    .Y(_2701_));
 sky130_fd_sc_hd__nor2_1 _6474_ (.A(_2701_),
    .B(_2700_),
    .Y(\egd_top.BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__nor2_1 _6475_ (.A(_3218_),
    .B(_3090_),
    .Y(_0182_));
 sky130_fd_sc_hd__xor2_2 _6476_ (.A(\egd_top.BitStream_buffer.pc_previous[4] ),
    .B(_2699_),
    .X(\egd_top.BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__nor2_1 _6477_ (.A(_3396_),
    .B(_3090_),
    .Y(_0181_));
 sky130_fd_sc_hd__nand2_2 _6478_ (.A(_2697_),
    .B(_2698_),
    .Y(_2702_));
 sky130_fd_sc_hd__xnor2_4 _6479_ (.A(_2702_),
    .B(_2696_),
    .Y(\egd_top.BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__nor2_1 _6480_ (.A(_3216_),
    .B(_3090_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_2 _6481_ (.A(_2694_),
    .B(_2695_),
    .Y(_2703_));
 sky130_fd_sc_hd__xnor2_4 _6482_ (.A(_2703_),
    .B(_2693_),
    .Y(\egd_top.BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__nor2_1 _6483_ (.A(_3276_),
    .B(_3090_),
    .Y(_0179_));
 sky130_fd_sc_hd__or2_1 _6484_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .X(_2704_));
 sky130_fd_sc_hd__and2_1 _6485_ (.A(_2704_),
    .B(_2692_),
    .X(_2705_));
 sky130_fd_sc_hd__xnor2_4 _6486_ (.A(_3113_),
    .B(_2705_),
    .Y(\egd_top.BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__nor2_1 _6487_ (.A(_3230_),
    .B(_3090_),
    .Y(_0178_));
 sky130_fd_sc_hd__nor2_1 _6488_ (.A(_3090_),
    .B(_3114_),
    .Y(_0177_));
 sky130_fd_sc_hd__nand3_4 _6489_ (.A(_3156_),
    .B(net42),
    .C(_2474_),
    .Y(_2706_));
 sky130_fd_sc_hd__clkbuf_4 _6490_ (.A(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__mux2_1 _6491_ (.A0(net7),
    .A1(_0781_),
    .S(_2707_),
    .X(_2708_));
 sky130_fd_sc_hd__and2_1 _6492_ (.A(_2708_),
    .B(_2689_),
    .X(_2709_));
 sky130_fd_sc_hd__clkbuf_1 _6493_ (.A(_2709_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _6494_ (.A0(net6),
    .A1(_0932_),
    .S(_2707_),
    .X(_2710_));
 sky130_fd_sc_hd__and2_1 _6495_ (.A(_2710_),
    .B(_2689_),
    .X(_2711_));
 sky130_fd_sc_hd__clkbuf_1 _6496_ (.A(_2711_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _6497_ (.A0(net5),
    .A1(_1073_),
    .S(_2707_),
    .X(_2712_));
 sky130_fd_sc_hd__and2_1 _6498_ (.A(_2712_),
    .B(_2689_),
    .X(_2713_));
 sky130_fd_sc_hd__clkbuf_1 _6499_ (.A(_2713_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _6500_ (.A0(net4),
    .A1(_1210_),
    .S(_2707_),
    .X(_2714_));
 sky130_fd_sc_hd__and2_1 _6501_ (.A(_2714_),
    .B(_2689_),
    .X(_2715_));
 sky130_fd_sc_hd__clkbuf_1 _6502_ (.A(_2715_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _6503_ (.A0(net3),
    .A1(_1055_),
    .S(_2707_),
    .X(_2716_));
 sky130_fd_sc_hd__and2_1 _6504_ (.A(_2716_),
    .B(_2689_),
    .X(_2717_));
 sky130_fd_sc_hd__clkbuf_1 _6505_ (.A(_2717_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _6506_ (.A0(net2),
    .A1(_1192_),
    .S(_2707_),
    .X(_2718_));
 sky130_fd_sc_hd__and2_1 _6507_ (.A(_2718_),
    .B(_2689_),
    .X(_2719_));
 sky130_fd_sc_hd__clkbuf_1 _6508_ (.A(_2719_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _6509_ (.A0(net16),
    .A1(_0510_),
    .S(_2707_),
    .X(_2720_));
 sky130_fd_sc_hd__and2_1 _6510_ (.A(_2720_),
    .B(_2689_),
    .X(_2721_));
 sky130_fd_sc_hd__clkbuf_1 _6511_ (.A(_2721_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _6512_ (.A0(net15),
    .A1(_0515_),
    .S(_2707_),
    .X(_2722_));
 sky130_fd_sc_hd__and2_1 _6513_ (.A(_2722_),
    .B(_2689_),
    .X(_2723_));
 sky130_fd_sc_hd__clkbuf_1 _6514_ (.A(_2723_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _6515_ (.A0(net14),
    .A1(_0765_),
    .S(_2707_),
    .X(_2724_));
 sky130_fd_sc_hd__and2_1 _6516_ (.A(_2724_),
    .B(_2689_),
    .X(_2725_));
 sky130_fd_sc_hd__clkbuf_1 _6517_ (.A(_2725_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _6518_ (.A0(net13),
    .A1(_0916_),
    .S(_2707_),
    .X(_2726_));
 sky130_fd_sc_hd__and2_1 _6519_ (.A(_2726_),
    .B(_3080_),
    .X(_2727_));
 sky130_fd_sc_hd__clkbuf_1 _6520_ (.A(_2727_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _6521_ (.A0(net12),
    .A1(_0518_),
    .S(_2706_),
    .X(_2728_));
 sky130_fd_sc_hd__and2_1 _6522_ (.A(_2728_),
    .B(_3080_),
    .X(_2729_));
 sky130_fd_sc_hd__clkbuf_1 _6523_ (.A(_2729_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(net11),
    .A1(_0522_),
    .S(_2706_),
    .X(_2730_));
 sky130_fd_sc_hd__and2_1 _6525_ (.A(_2730_),
    .B(_3080_),
    .X(_2731_));
 sky130_fd_sc_hd__clkbuf_1 _6526_ (.A(_2731_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _6527_ (.A0(net10),
    .A1(_0768_),
    .S(_2706_),
    .X(_2732_));
 sky130_fd_sc_hd__and2_1 _6528_ (.A(_2732_),
    .B(_3080_),
    .X(_2733_));
 sky130_fd_sc_hd__clkbuf_1 _6529_ (.A(_2733_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _6530_ (.A0(net9),
    .A1(_0919_),
    .S(_2706_),
    .X(_2734_));
 sky130_fd_sc_hd__and2_1 _6531_ (.A(_2734_),
    .B(_3080_),
    .X(_2735_));
 sky130_fd_sc_hd__clkbuf_1 _6532_ (.A(_2735_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _6533_ (.A0(net8),
    .A1(_0534_),
    .S(_2706_),
    .X(_2736_));
 sky130_fd_sc_hd__and2_1 _6534_ (.A(_2736_),
    .B(_3080_),
    .X(_2737_));
 sky130_fd_sc_hd__clkbuf_1 _6535_ (.A(_2737_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _6536_ (.A0(net1),
    .A1(_0538_),
    .S(_2706_),
    .X(_2738_));
 sky130_fd_sc_hd__and2_1 _6537_ (.A(_2738_),
    .B(_3080_),
    .X(_2739_));
 sky130_fd_sc_hd__clkbuf_1 _6538_ (.A(_2739_),
    .X(_0161_));
 sky130_fd_sc_hd__inv_2 _6539_ (.A(_3111_),
    .Y(_2740_));
 sky130_fd_sc_hd__nand2_1 _6540_ (.A(net18),
    .B(net17),
    .Y(_2741_));
 sky130_fd_sc_hd__inv_2 _6541_ (.A(_2741_),
    .Y(_2742_));
 sky130_fd_sc_hd__and3b_1 _6542_ (.A_N(net25),
    .B(_2742_),
    .C(net24),
    .X(_2743_));
 sky130_fd_sc_hd__inv_2 _6543_ (.A(\egd_top.exp_golomb_decoding.te_range[2] ),
    .Y(_2744_));
 sky130_fd_sc_hd__and2_1 _6544_ (.A(_2743_),
    .B(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__inv_2 _6545_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2746_));
 sky130_fd_sc_hd__nand2_1 _6546_ (.A(_2746_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2747_));
 sky130_fd_sc_hd__inv_2 _6547_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2748_));
 sky130_fd_sc_hd__nand2_1 _6548_ (.A(_2747_),
    .B(_2748_),
    .Y(_2749_));
 sky130_fd_sc_hd__inv_2 _6549_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2750_));
 sky130_fd_sc_hd__nand2_1 _6550_ (.A(_2749_),
    .B(_2750_),
    .Y(_2751_));
 sky130_fd_sc_hd__inv_2 _6551_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2752_));
 sky130_fd_sc_hd__nand2_1 _6552_ (.A(_2751_),
    .B(_2752_),
    .Y(_2753_));
 sky130_fd_sc_hd__inv_2 _6553_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2754_));
 sky130_fd_sc_hd__nand2_1 _6554_ (.A(_2753_),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__inv_2 _6555_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2756_));
 sky130_fd_sc_hd__nand2_1 _6556_ (.A(_2755_),
    .B(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__inv_2 _6557_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_2758_));
 sky130_fd_sc_hd__nand2_1 _6558_ (.A(_2757_),
    .B(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__inv_2 _6559_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2760_));
 sky130_fd_sc_hd__nand2_1 _6560_ (.A(_2759_),
    .B(_2760_),
    .Y(_2761_));
 sky130_fd_sc_hd__inv_2 _6561_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2762_));
 sky130_fd_sc_hd__inv_4 _6562_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2763_));
 sky130_fd_sc_hd__nand2_1 _6563_ (.A(_2762_),
    .B(_2763_),
    .Y(_2764_));
 sky130_fd_sc_hd__nor2_1 _6564_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__inv_2 _6565_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_2766_));
 sky130_fd_sc_hd__nand2_2 _6566_ (.A(_2765_),
    .B(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hd__inv_2 _6567_ (.A(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__nand2_1 _6568_ (.A(_2761_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__a21oi_1 _6569_ (.A1(_2762_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2770_));
 sky130_fd_sc_hd__nand2_1 _6570_ (.A(_2769_),
    .B(_2770_),
    .Y(_2771_));
 sky130_fd_sc_hd__nor2_1 _6571_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2772_));
 sky130_fd_sc_hd__nand2_2 _6572_ (.A(_2771_),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__nor2_1 _6573_ (.A(_3149_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_2774_));
 sky130_fd_sc_hd__nand2_1 _6574_ (.A(_2773_),
    .B(_2774_),
    .Y(_2775_));
 sky130_fd_sc_hd__or3_1 _6575_ (.A(_2740_),
    .B(_2745_),
    .C(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__inv_2 _6576_ (.A(_2776_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__o21a_1 _6577_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_2750_),
    .X(_2777_));
 sky130_fd_sc_hd__a211o_1 _6578_ (.A1(_2777_),
    .A2(_2752_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .C1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .X(_2778_));
 sky130_fd_sc_hd__and3_2 _6579_ (.A(_2768_),
    .B(_2760_),
    .C(_2758_),
    .X(_2779_));
 sky130_fd_sc_hd__nor2_2 _6580_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2780_));
 sky130_fd_sc_hd__nand2_1 _6581_ (.A(_2772_),
    .B(_3150_),
    .Y(_2781_));
 sky130_fd_sc_hd__a21o_1 _6582_ (.A1(_2767_),
    .A2(_2780_),
    .B1(_2781_),
    .X(_2782_));
 sky130_fd_sc_hd__a21oi_4 _6583_ (.A1(_2778_),
    .A2(_2779_),
    .B1(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__clkinvlp_2 _6584_ (.A(_2783_),
    .Y(_2784_));
 sky130_fd_sc_hd__or3_1 _6585_ (.A(_2740_),
    .B(_2745_),
    .C(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__inv_2 _6586_ (.A(_2785_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__nor2_1 _6587_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2786_));
 sky130_fd_sc_hd__inv_2 _6588_ (.A(_2786_),
    .Y(_2787_));
 sky130_fd_sc_hd__nor2_1 _6589_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__nand2_1 _6590_ (.A(_2788_),
    .B(_2750_),
    .Y(_2789_));
 sky130_fd_sc_hd__nand2_1 _6591_ (.A(_2779_),
    .B(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__inv_2 _6592_ (.A(_2781_),
    .Y(_2791_));
 sky130_fd_sc_hd__nand2_1 _6593_ (.A(_2791_),
    .B(_2780_),
    .Y(_2792_));
 sky130_fd_sc_hd__inv_2 _6594_ (.A(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__nand2_1 _6595_ (.A(_2790_),
    .B(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__or3_1 _6596_ (.A(_2740_),
    .B(_2745_),
    .C(_2794_),
    .X(_2795_));
 sky130_fd_sc_hd__inv_2 _6597_ (.A(_2795_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__nand2_1 _6598_ (.A(_2760_),
    .B(_2758_),
    .Y(_2796_));
 sky130_fd_sc_hd__o211ai_4 _6599_ (.A1(_2796_),
    .A2(_2767_),
    .B1(_2780_),
    .C1(_2791_),
    .Y(_2797_));
 sky130_fd_sc_hd__or2_1 _6600_ (.A(_2783_),
    .B(_2775_),
    .X(_2798_));
 sky130_fd_sc_hd__nor2_2 _6601_ (.A(_2797_),
    .B(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__nor2_1 _6602_ (.A(_2797_),
    .B(_2783_),
    .Y(_2800_));
 sky130_fd_sc_hd__nand2_2 _6603_ (.A(_2775_),
    .B(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__nand2_1 _6604_ (.A(_2783_),
    .B(_2792_),
    .Y(_2802_));
 sky130_fd_sc_hd__a21oi_1 _6605_ (.A1(_2773_),
    .A2(_2774_),
    .B1(_2802_),
    .Y(_2803_));
 sky130_fd_sc_hd__nand2_1 _6606_ (.A(_2803_),
    .B(_2763_),
    .Y(_2804_));
 sky130_fd_sc_hd__o21ai_1 _6607_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .A2(_2801_),
    .B1(_2804_),
    .Y(_2805_));
 sky130_fd_sc_hd__a21oi_1 _6608_ (.A1(_2799_),
    .A2(_2752_),
    .B1(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__nor2_1 _6609_ (.A(_2793_),
    .B(_2798_),
    .Y(_2807_));
 sky130_fd_sc_hd__inv_2 _6610_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2808_));
 sky130_fd_sc_hd__nand3_4 _6611_ (.A(_2773_),
    .B(_2774_),
    .C(_2783_),
    .Y(_2809_));
 sky130_fd_sc_hd__nor2_1 _6612_ (.A(_2793_),
    .B(_2809_),
    .Y(_2810_));
 sky130_fd_sc_hd__and2_1 _6613_ (.A(_2810_),
    .B(_2760_),
    .X(_2811_));
 sky130_fd_sc_hd__a21oi_1 _6614_ (.A1(_2807_),
    .A2(_2808_),
    .B1(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__o21ai_1 _6615_ (.A1(_2797_),
    .A2(_2809_),
    .B1(_2748_),
    .Y(_2813_));
 sky130_fd_sc_hd__nor2_4 _6616_ (.A(_2797_),
    .B(_2809_),
    .Y(_2814_));
 sky130_fd_sc_hd__inv_2 _6617_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2815_));
 sky130_fd_sc_hd__nand2_1 _6618_ (.A(_2814_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__nand2_2 _6619_ (.A(_2813_),
    .B(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__nor2_2 _6620_ (.A(_2797_),
    .B(_2784_),
    .Y(_2818_));
 sky130_fd_sc_hd__nand2_1 _6621_ (.A(_2817_),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__nand3_2 _6622_ (.A(_2806_),
    .B(_2812_),
    .C(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__inv_2 _6623_ (.A(_2779_),
    .Y(_2821_));
 sky130_fd_sc_hd__nor2_1 _6624_ (.A(_2781_),
    .B(_2821_),
    .Y(_2822_));
 sky130_fd_sc_hd__and3_1 _6625_ (.A(_2775_),
    .B(_2784_),
    .C(_2794_),
    .X(_2823_));
 sky130_fd_sc_hd__or3_1 _6626_ (.A(_2740_),
    .B(_2822_),
    .C(_2823_),
    .X(_2824_));
 sky130_fd_sc_hd__inv_2 _6627_ (.A(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__o211a_1 _6628_ (.A1(_2745_),
    .A2(_2820_),
    .B1(_2742_),
    .C1(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__o21ai_1 _6629_ (.A1(_2797_),
    .A2(_2809_),
    .B1(_2750_),
    .Y(_2827_));
 sky130_fd_sc_hd__inv_2 _6630_ (.A(_2809_),
    .Y(_2828_));
 sky130_fd_sc_hd__inv_2 _6631_ (.A(_2797_),
    .Y(_2829_));
 sky130_fd_sc_hd__nand3_1 _6632_ (.A(_2828_),
    .B(_2746_),
    .C(_2829_),
    .Y(_2830_));
 sky130_fd_sc_hd__nand2_2 _6633_ (.A(_2827_),
    .B(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__nand3_1 _6634_ (.A(_2831_),
    .B(_2813_),
    .C(_2816_),
    .Y(_2832_));
 sky130_fd_sc_hd__nand2_2 _6635_ (.A(_2828_),
    .B(_2829_),
    .Y(_2833_));
 sky130_fd_sc_hd__nand2_1 _6636_ (.A(_2833_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2834_));
 sky130_fd_sc_hd__nand2_1 _6637_ (.A(_2814_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2835_));
 sky130_fd_sc_hd__nand2_1 _6638_ (.A(_2834_),
    .B(_2835_),
    .Y(_2836_));
 sky130_fd_sc_hd__nand2_1 _6639_ (.A(_2836_),
    .B(_2817_),
    .Y(_2837_));
 sky130_fd_sc_hd__nand3_1 _6640_ (.A(_2832_),
    .B(_2837_),
    .C(_2818_),
    .Y(_2838_));
 sky130_fd_sc_hd__xnor2_1 _6641_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2839_));
 sky130_fd_sc_hd__nand2_1 _6642_ (.A(_2807_),
    .B(_2839_),
    .Y(_2840_));
 sky130_fd_sc_hd__nor2_1 _6643_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2841_));
 sky130_fd_sc_hd__inv_2 _6644_ (.A(_2841_),
    .Y(_2842_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2843_));
 sky130_fd_sc_hd__nand2_1 _6646_ (.A(_2842_),
    .B(_2843_),
    .Y(_2844_));
 sky130_fd_sc_hd__nand2_1 _6647_ (.A(_2810_),
    .B(_2844_),
    .Y(_2845_));
 sky130_fd_sc_hd__nand2_1 _6648_ (.A(_2840_),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__nor2_1 _6649_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2847_));
 sky130_fd_sc_hd__inv_2 _6650_ (.A(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__nand2_1 _6651_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2849_));
 sky130_fd_sc_hd__and2_1 _6652_ (.A(_2848_),
    .B(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__xnor2_1 _6653_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2851_));
 sky130_fd_sc_hd__nand2_1 _6654_ (.A(_2803_),
    .B(_2851_),
    .Y(_2852_));
 sky130_fd_sc_hd__o21ai_1 _6655_ (.A1(_2801_),
    .A2(_2850_),
    .B1(_2852_),
    .Y(_2853_));
 sky130_fd_sc_hd__inv_2 _6656_ (.A(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__nand2_1 _6657_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2855_));
 sky130_fd_sc_hd__nand2_1 _6658_ (.A(_2787_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__nand2_1 _6659_ (.A(_2799_),
    .B(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__nand2_1 _6660_ (.A(_2854_),
    .B(_2857_),
    .Y(_2858_));
 sky130_fd_sc_hd__nor2_1 _6661_ (.A(_2846_),
    .B(_2858_),
    .Y(_2859_));
 sky130_fd_sc_hd__nand2_1 _6662_ (.A(_2838_),
    .B(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__buf_2 _6663_ (.A(_3111_),
    .X(_2861_));
 sky130_fd_sc_hd__nand3_1 _6664_ (.A(_2860_),
    .B(_2861_),
    .C(_2820_),
    .Y(_2862_));
 sky130_fd_sc_hd__inv_2 _6665_ (.A(_2862_),
    .Y(_2863_));
 sky130_fd_sc_hd__nand2_2 _6666_ (.A(_2820_),
    .B(_2861_),
    .Y(_2864_));
 sky130_fd_sc_hd__inv_4 _6667_ (.A(_2864_),
    .Y(_2865_));
 sky130_fd_sc_hd__nand2_1 _6668_ (.A(_2860_),
    .B(_2861_),
    .Y(_2866_));
 sky130_fd_sc_hd__inv_2 _6669_ (.A(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__nor2_1 _6670_ (.A(_2865_),
    .B(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__nor2_2 _6671_ (.A(net17),
    .B(_3109_),
    .Y(_2869_));
 sky130_fd_sc_hd__or3b_1 _6672_ (.A(_2863_),
    .B(_2868_),
    .C_N(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__or3_1 _6673_ (.A(net18),
    .B(_3110_),
    .C(_2864_),
    .X(_2871_));
 sky130_fd_sc_hd__nand3b_2 _6674_ (.A_N(_2826_),
    .B(_2870_),
    .C(_2871_),
    .Y(net24));
 sky130_fd_sc_hd__nand2_2 _6675_ (.A(_2817_),
    .B(_2831_),
    .Y(_2872_));
 sky130_fd_sc_hd__nand2_1 _6676_ (.A(_2833_),
    .B(_2752_),
    .Y(_2873_));
 sky130_fd_sc_hd__nand2_1 _6677_ (.A(_2814_),
    .B(_2748_),
    .Y(_2874_));
 sky130_fd_sc_hd__nand2_1 _6678_ (.A(_2873_),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__nand2_1 _6679_ (.A(_2872_),
    .B(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__o21ai_1 _6680_ (.A1(_2797_),
    .A2(_2809_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2877_));
 sky130_fd_sc_hd__nand2_1 _6681_ (.A(_2814_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2878_));
 sky130_fd_sc_hd__nand2_1 _6682_ (.A(_2877_),
    .B(_2878_),
    .Y(_2879_));
 sky130_fd_sc_hd__nand3_1 _6683_ (.A(_2817_),
    .B(_2879_),
    .C(_2831_),
    .Y(_2880_));
 sky130_fd_sc_hd__nand3_1 _6684_ (.A(_2876_),
    .B(_2880_),
    .C(_2818_),
    .Y(_2881_));
 sky130_fd_sc_hd__nand2_1 _6685_ (.A(_2847_),
    .B(_2760_),
    .Y(_2882_));
 sky130_fd_sc_hd__nand2_1 _6686_ (.A(_2848_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2883_));
 sky130_fd_sc_hd__a21o_1 _6687_ (.A1(_2882_),
    .A2(_2883_),
    .B1(_2801_),
    .X(_2884_));
 sky130_fd_sc_hd__and2_1 _6688_ (.A(_2764_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .X(_2885_));
 sky130_fd_sc_hd__o21ai_1 _6689_ (.A1(_2765_),
    .A2(_2885_),
    .B1(_2803_),
    .Y(_2886_));
 sky130_fd_sc_hd__nand2_1 _6690_ (.A(_2884_),
    .B(_2886_),
    .Y(_2887_));
 sky130_fd_sc_hd__nor2_1 _6691_ (.A(_2756_),
    .B(_2786_),
    .Y(_2888_));
 sky130_fd_sc_hd__o21ai_1 _6692_ (.A1(_2788_),
    .A2(_2888_),
    .B1(_2799_),
    .Y(_2889_));
 sky130_fd_sc_hd__nor2_1 _6693_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2842_),
    .Y(_2890_));
 sky130_fd_sc_hd__nor2_1 _6694_ (.A(_2763_),
    .B(_2841_),
    .Y(_2891_));
 sky130_fd_sc_hd__o21ai_1 _6695_ (.A1(_2890_),
    .A2(_2891_),
    .B1(_2810_),
    .Y(_2892_));
 sky130_fd_sc_hd__nand2_1 _6696_ (.A(_2889_),
    .B(_2892_),
    .Y(_2893_));
 sky130_fd_sc_hd__nor2_1 _6697_ (.A(_2887_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__nand2_1 _6698_ (.A(_2881_),
    .B(_2894_),
    .Y(_2895_));
 sky130_fd_sc_hd__o21ai_1 _6699_ (.A1(_2860_),
    .A2(_2895_),
    .B1(_2861_),
    .Y(_2896_));
 sky130_fd_sc_hd__inv_2 _6700_ (.A(_2896_),
    .Y(_2897_));
 sky130_fd_sc_hd__nand3_1 _6701_ (.A(_2895_),
    .B(_2861_),
    .C(_2860_),
    .Y(_2898_));
 sky130_fd_sc_hd__a31o_1 _6702_ (.A1(_2743_),
    .A2(net18),
    .A3(_2744_),
    .B1(_3110_),
    .X(_2899_));
 sky130_fd_sc_hd__inv_2 _6703_ (.A(_2899_),
    .Y(_2900_));
 sky130_fd_sc_hd__a32o_2 _6704_ (.A1(_2897_),
    .A2(_2898_),
    .A3(_2869_),
    .B1(_2867_),
    .B2(_2900_),
    .X(net25));
 sky130_fd_sc_hd__nand2_1 _6705_ (.A(_2898_),
    .B(_2865_),
    .Y(_2901_));
 sky130_fd_sc_hd__nand2_1 _6706_ (.A(_2897_),
    .B(_2901_),
    .Y(_2902_));
 sky130_fd_sc_hd__inv_2 _6707_ (.A(_2872_),
    .Y(_2903_));
 sky130_fd_sc_hd__nand2_1 _6708_ (.A(_2833_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2904_));
 sky130_fd_sc_hd__nand2_1 _6709_ (.A(_2814_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2905_));
 sky130_fd_sc_hd__nand2_1 _6710_ (.A(_2904_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__nand3_1 _6711_ (.A(_2903_),
    .B(_2875_),
    .C(_2906_),
    .Y(_2907_));
 sky130_fd_sc_hd__nand3_1 _6712_ (.A(_2875_),
    .B(_2817_),
    .C(_2831_),
    .Y(_2908_));
 sky130_fd_sc_hd__o21ai_1 _6713_ (.A1(_2797_),
    .A2(_2809_),
    .B1(_2754_),
    .Y(_2909_));
 sky130_fd_sc_hd__nand2_1 _6714_ (.A(_2814_),
    .B(_2750_),
    .Y(_2910_));
 sky130_fd_sc_hd__nand2_1 _6715_ (.A(_2909_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__nand2_1 _6716_ (.A(_2908_),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__nand3_1 _6717_ (.A(_2907_),
    .B(_2818_),
    .C(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__nor2_1 _6718_ (.A(_2787_),
    .B(_2848_),
    .Y(_2914_));
 sky130_fd_sc_hd__nor2_1 _6719_ (.A(_2758_),
    .B(_2788_),
    .Y(_2915_));
 sky130_fd_sc_hd__o21ai_1 _6720_ (.A1(_2914_),
    .A2(_2915_),
    .B1(_2799_),
    .Y(_2916_));
 sky130_fd_sc_hd__nand2_1 _6721_ (.A(_2890_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2917_));
 sky130_fd_sc_hd__or2_1 _6722_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(_2890_),
    .X(_2918_));
 sky130_fd_sc_hd__nand3_1 _6723_ (.A(_2810_),
    .B(_2917_),
    .C(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__nand2_1 _6724_ (.A(_2847_),
    .B(_2841_),
    .Y(_2920_));
 sky130_fd_sc_hd__nand2_1 _6725_ (.A(_2882_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_2921_));
 sky130_fd_sc_hd__a21o_1 _6726_ (.A1(_2920_),
    .A2(_2921_),
    .B1(_2801_),
    .X(_2922_));
 sky130_fd_sc_hd__and3_1 _6727_ (.A(_2916_),
    .B(_2919_),
    .C(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__a21oi_1 _6728_ (.A1(_2913_),
    .A2(_2923_),
    .B1(_2740_),
    .Y(_2924_));
 sky130_fd_sc_hd__nand2_1 _6729_ (.A(_2902_),
    .B(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__nand2_1 _6730_ (.A(_2913_),
    .B(_2923_),
    .Y(_2926_));
 sky130_fd_sc_hd__nand2_1 _6731_ (.A(_2926_),
    .B(_2861_),
    .Y(_2927_));
 sky130_fd_sc_hd__nand3_1 _6732_ (.A(_2897_),
    .B(_2927_),
    .C(_2901_),
    .Y(_2928_));
 sky130_fd_sc_hd__nand2_1 _6733_ (.A(_2925_),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__nand2_1 _6734_ (.A(_2929_),
    .B(_2869_),
    .Y(_2930_));
 sky130_fd_sc_hd__nand2_1 _6735_ (.A(_2895_),
    .B(_2861_),
    .Y(_2931_));
 sky130_fd_sc_hd__inv_2 _6736_ (.A(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__nand2_1 _6737_ (.A(_2932_),
    .B(_2900_),
    .Y(_2933_));
 sky130_fd_sc_hd__nand2_1 _6738_ (.A(net24),
    .B(net25),
    .Y(_2934_));
 sky130_fd_sc_hd__a21oi_1 _6739_ (.A1(_2930_),
    .A2(_2933_),
    .B1(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__nand3_1 _6740_ (.A(_2930_),
    .B(_2934_),
    .C(_2933_),
    .Y(_2936_));
 sky130_fd_sc_hd__nand2_1 _6741_ (.A(_2936_),
    .B(_2742_),
    .Y(_2937_));
 sky130_fd_sc_hd__nor2_1 _6742_ (.A(_2935_),
    .B(_2937_),
    .Y(\egd_top.exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__nand2_1 _6743_ (.A(_2930_),
    .B(_2933_),
    .Y(net26));
 sky130_fd_sc_hd__nand2_1 _6744_ (.A(_2875_),
    .B(_2911_),
    .Y(_2938_));
 sky130_fd_sc_hd__nand2_1 _6745_ (.A(_2814_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2939_));
 sky130_fd_sc_hd__o21ai_2 _6746_ (.A1(_2756_),
    .A2(_2814_),
    .B1(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__inv_2 _6747_ (.A(_2940_),
    .Y(_2941_));
 sky130_fd_sc_hd__o21ai_1 _6748_ (.A1(_2872_),
    .A2(_2938_),
    .B1(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__nor2_1 _6749_ (.A(_2872_),
    .B(_2938_),
    .Y(_2943_));
 sky130_fd_sc_hd__nand2_1 _6750_ (.A(_2943_),
    .B(_2940_),
    .Y(_2944_));
 sky130_fd_sc_hd__nand3_1 _6751_ (.A(_2942_),
    .B(_2944_),
    .C(_2818_),
    .Y(_2945_));
 sky130_fd_sc_hd__and2_1 _6752_ (.A(_2920_),
    .B(_2763_),
    .X(_2946_));
 sky130_fd_sc_hd__nor2_1 _6753_ (.A(_2763_),
    .B(_2920_),
    .Y(_2947_));
 sky130_fd_sc_hd__nor2_1 _6754_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2914_),
    .Y(_2948_));
 sky130_fd_sc_hd__inv_2 _6755_ (.A(_2914_),
    .Y(_2949_));
 sky130_fd_sc_hd__nor2_1 _6756_ (.A(_2760_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__or2_1 _6757_ (.A(_2948_),
    .B(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__inv_2 _6758_ (.A(_2799_),
    .Y(_2952_));
 sky130_fd_sc_hd__o32a_1 _6759_ (.A1(_2946_),
    .A2(_2801_),
    .A3(_2947_),
    .B1(_2951_),
    .B2(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__a21oi_2 _6760_ (.A1(_2945_),
    .A2(_2953_),
    .B1(_2740_),
    .Y(_2954_));
 sky130_fd_sc_hd__inv_2 _6761_ (.A(_2954_),
    .Y(_2955_));
 sky130_fd_sc_hd__nand2_1 _6762_ (.A(_2896_),
    .B(_2927_),
    .Y(_2956_));
 sky130_fd_sc_hd__nor2_1 _6763_ (.A(_2931_),
    .B(_2862_),
    .Y(_2957_));
 sky130_fd_sc_hd__nand2_1 _6764_ (.A(_2924_),
    .B(_2957_),
    .Y(_2958_));
 sky130_fd_sc_hd__nand2_1 _6765_ (.A(_2958_),
    .B(_2865_),
    .Y(_2959_));
 sky130_fd_sc_hd__o21ai_1 _6766_ (.A1(_2865_),
    .A2(_2956_),
    .B1(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__or2_1 _6767_ (.A(_2955_),
    .B(_2960_),
    .X(_2961_));
 sky130_fd_sc_hd__nand2_1 _6768_ (.A(_2960_),
    .B(_2955_),
    .Y(_2962_));
 sky130_fd_sc_hd__nand3_1 _6769_ (.A(_2961_),
    .B(_2869_),
    .C(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__nand2_1 _6770_ (.A(_2924_),
    .B(_2900_),
    .Y(_2964_));
 sky130_fd_sc_hd__nand2_1 _6771_ (.A(_2963_),
    .B(_2964_),
    .Y(net27));
 sky130_fd_sc_hd__o21ai_1 _6772_ (.A1(_2958_),
    .A2(_2955_),
    .B1(_2865_),
    .Y(_2965_));
 sky130_fd_sc_hd__nor2_1 _6773_ (.A(_2954_),
    .B(_2956_),
    .Y(_2966_));
 sky130_fd_sc_hd__nand2_1 _6774_ (.A(_2966_),
    .B(_2864_),
    .Y(_2967_));
 sky130_fd_sc_hd__nand2_1 _6775_ (.A(_2965_),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__nor2_1 _6776_ (.A(_2879_),
    .B(_2906_),
    .Y(_2969_));
 sky130_fd_sc_hd__nand3_1 _6777_ (.A(_2903_),
    .B(_2969_),
    .C(_2941_),
    .Y(_2970_));
 sky130_fd_sc_hd__a21oi_2 _6778_ (.A1(_2814_),
    .A2(_2754_),
    .B1(_2758_),
    .Y(_2971_));
 sky130_fd_sc_hd__inv_2 _6779_ (.A(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__nand2_1 _6780_ (.A(_2970_),
    .B(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__nand3_1 _6781_ (.A(_2943_),
    .B(_2941_),
    .C(_2971_),
    .Y(_2974_));
 sky130_fd_sc_hd__nand3_1 _6782_ (.A(_2973_),
    .B(_2974_),
    .C(_2818_),
    .Y(_2975_));
 sky130_fd_sc_hd__nor2_1 _6783_ (.A(_2844_),
    .B(_2949_),
    .Y(_2976_));
 sky130_fd_sc_hd__a211o_1 _6784_ (.A1(_2766_),
    .A2(_2949_),
    .B1(_2976_),
    .C1(_2952_),
    .X(_2977_));
 sky130_fd_sc_hd__nand2_1 _6785_ (.A(_2975_),
    .B(_2977_),
    .Y(_2978_));
 sky130_fd_sc_hd__nand2_1 _6786_ (.A(_2978_),
    .B(_2861_),
    .Y(_2979_));
 sky130_fd_sc_hd__nand2_1 _6787_ (.A(_2968_),
    .B(_2979_),
    .Y(_2980_));
 sky130_fd_sc_hd__inv_2 _6788_ (.A(_2979_),
    .Y(_2981_));
 sky130_fd_sc_hd__nand3_1 _6789_ (.A(_2965_),
    .B(_2981_),
    .C(_2967_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand3_1 _6790_ (.A(_2980_),
    .B(_2869_),
    .C(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__nand2_1 _6791_ (.A(_2954_),
    .B(_2900_),
    .Y(_2984_));
 sky130_fd_sc_hd__nand2_1 _6792_ (.A(_2983_),
    .B(_2984_),
    .Y(net28));
 sky130_fd_sc_hd__nand2_1 _6793_ (.A(_2945_),
    .B(_2953_),
    .Y(_2985_));
 sky130_fd_sc_hd__nand3_1 _6794_ (.A(_2978_),
    .B(_2861_),
    .C(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__o21ai_1 _6795_ (.A1(_2958_),
    .A2(_2986_),
    .B1(_2865_),
    .Y(_2987_));
 sky130_fd_sc_hd__nand3_1 _6796_ (.A(_2966_),
    .B(_2864_),
    .C(_2979_),
    .Y(_2988_));
 sky130_fd_sc_hd__nand2_1 _6797_ (.A(_2987_),
    .B(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__inv_2 _6798_ (.A(_2818_),
    .Y(_2990_));
 sky130_fd_sc_hd__nor2_1 _6799_ (.A(_2971_),
    .B(_2940_),
    .Y(_2991_));
 sky130_fd_sc_hd__nand2_1 _6800_ (.A(_2943_),
    .B(_2991_),
    .Y(_2992_));
 sky130_fd_sc_hd__o21ai_2 _6801_ (.A1(_2756_),
    .A2(_2833_),
    .B1(_2760_),
    .Y(_2993_));
 sky130_fd_sc_hd__inv_2 _6802_ (.A(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__nand2_1 _6803_ (.A(_2992_),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__nand3_1 _6804_ (.A(_2943_),
    .B(_2991_),
    .C(_2993_),
    .Y(_2996_));
 sky130_fd_sc_hd__nand2_1 _6805_ (.A(_2995_),
    .B(_2996_),
    .Y(_2997_));
 sky130_fd_sc_hd__nor2_1 _6806_ (.A(_2990_),
    .B(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__and2_1 _6807_ (.A(_2998_),
    .B(_2825_),
    .X(_2999_));
 sky130_fd_sc_hd__inv_2 _6808_ (.A(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__nand2_1 _6809_ (.A(_2989_),
    .B(_3000_),
    .Y(_3001_));
 sky130_fd_sc_hd__nand3_1 _6810_ (.A(_2987_),
    .B(_2988_),
    .C(_2999_),
    .Y(_3002_));
 sky130_fd_sc_hd__nand3_1 _6811_ (.A(_3001_),
    .B(_3002_),
    .C(_2869_),
    .Y(_3003_));
 sky130_fd_sc_hd__nand2_1 _6812_ (.A(_2981_),
    .B(_2900_),
    .Y(_3004_));
 sky130_fd_sc_hd__nand2_1 _6813_ (.A(_3003_),
    .B(_3004_),
    .Y(net29));
 sky130_fd_sc_hd__inv_2 _6814_ (.A(_2986_),
    .Y(_3005_));
 sky130_fd_sc_hd__nand2_1 _6815_ (.A(_2863_),
    .B(_2932_),
    .Y(_3006_));
 sky130_fd_sc_hd__nor2_1 _6816_ (.A(_2927_),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__nand3_1 _6817_ (.A(_3005_),
    .B(_2999_),
    .C(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__o21ai_1 _6818_ (.A1(_2993_),
    .A2(_2992_),
    .B1(_2814_),
    .Y(_3009_));
 sky130_fd_sc_hd__inv_2 _6819_ (.A(_3009_),
    .Y(_3010_));
 sky130_fd_sc_hd__nand2_1 _6820_ (.A(_3010_),
    .B(_2825_),
    .Y(_3011_));
 sky130_fd_sc_hd__nand2_1 _6821_ (.A(_3008_),
    .B(_3011_),
    .Y(_3012_));
 sky130_fd_sc_hd__nand2_1 _6822_ (.A(_3012_),
    .B(_2865_),
    .Y(_3013_));
 sky130_fd_sc_hd__o21ai_1 _6823_ (.A1(_2998_),
    .A2(_2978_),
    .B1(_2861_),
    .Y(_3014_));
 sky130_fd_sc_hd__nand2_1 _6824_ (.A(_3014_),
    .B(_2966_),
    .Y(_3015_));
 sky130_fd_sc_hd__inv_2 _6825_ (.A(_3011_),
    .Y(_3016_));
 sky130_fd_sc_hd__nand2_1 _6826_ (.A(_3015_),
    .B(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__nor2_1 _6827_ (.A(_2824_),
    .B(_2820_),
    .Y(_3018_));
 sky130_fd_sc_hd__nand2_1 _6828_ (.A(_3017_),
    .B(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__nand2_1 _6829_ (.A(_3013_),
    .B(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__nand2_1 _6830_ (.A(_3020_),
    .B(_2869_),
    .Y(_3021_));
 sky130_fd_sc_hd__nand2_1 _6831_ (.A(_2999_),
    .B(_2900_),
    .Y(_3022_));
 sky130_fd_sc_hd__nand2_1 _6832_ (.A(_3021_),
    .B(_3022_),
    .Y(net30));
 sky130_fd_sc_hd__a22o_1 _6833_ (.A1(_2869_),
    .A2(_3018_),
    .B1(_3016_),
    .B2(_2900_),
    .X(net31));
 sky130_fd_sc_hd__buf_4 _6834_ (.A(net19),
    .X(_3023_));
 sky130_fd_sc_hd__clkbuf_8 _6835_ (.A(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__buf_4 _6836_ (.A(_3024_),
    .X(_3025_));
 sky130_fd_sc_hd__clkbuf_8 _6837_ (.A(net21),
    .X(_3026_));
 sky130_fd_sc_hd__buf_4 _6838_ (.A(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__buf_4 _6839_ (.A(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__or2b_2 _6840_ (.A(wb_clk_i),
    .B_N(_3026_),
    .X(_3029_));
 sky130_fd_sc_hd__buf_1 _6841_ (.A(_3029_),
    .X(_3030_));
 sky130_fd_sc_hd__buf_1 _6842_ (.A(clknet_1_1__leaf__3030_),
    .X(_3031_));
 sky130_fd_sc_hd__buf_1 _6843_ (.A(clknet_1_0__leaf__3031_),
    .X(_3032_));
 sky130_fd_sc_hd__o21ai_2 _6844_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_1__leaf__3032_),
    .Y(_0000_));
 sky130_fd_sc_hd__o21ai_2 _6845_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_1__leaf__3032_),
    .Y(_0001_));
 sky130_fd_sc_hd__o21ai_2 _6846_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_1__leaf__3032_),
    .Y(_0002_));
 sky130_fd_sc_hd__o21ai_2 _6847_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_1__leaf__3032_),
    .Y(_0003_));
 sky130_fd_sc_hd__o21ai_2 _6848_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_1__leaf__3032_),
    .Y(_0004_));
 sky130_fd_sc_hd__o21ai_2 _6849_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_0__leaf__3032_),
    .Y(_0005_));
 sky130_fd_sc_hd__o21ai_2 _6850_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_0__leaf__3032_),
    .Y(_0006_));
 sky130_fd_sc_hd__o21ai_2 _6851_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_0__leaf__3032_),
    .Y(_0007_));
 sky130_fd_sc_hd__o21ai_2 _6852_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_0__leaf__3032_),
    .Y(_0008_));
 sky130_fd_sc_hd__o21ai_2 _6853_ (.A1(_3025_),
    .A2(_3028_),
    .B1(clknet_1_0__leaf__3032_),
    .Y(_0009_));
 sky130_fd_sc_hd__buf_4 _6854_ (.A(_3024_),
    .X(_3033_));
 sky130_fd_sc_hd__buf_4 _6855_ (.A(_3027_),
    .X(_3034_));
 sky130_fd_sc_hd__buf_1 _6856_ (.A(clknet_1_0__leaf__3031_),
    .X(_3035_));
 sky130_fd_sc_hd__o21ai_2 _6857_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_0__leaf__3035_),
    .Y(_0010_));
 sky130_fd_sc_hd__o21ai_2 _6858_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_0__leaf__3035_),
    .Y(_0011_));
 sky130_fd_sc_hd__o21ai_2 _6859_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_0__leaf__3035_),
    .Y(_0012_));
 sky130_fd_sc_hd__o21ai_2 _6860_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_1__leaf__3035_),
    .Y(_0013_));
 sky130_fd_sc_hd__o21ai_2 _6861_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_1__leaf__3035_),
    .Y(_0014_));
 sky130_fd_sc_hd__o21ai_2 _6862_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_1__leaf__3035_),
    .Y(_0015_));
 sky130_fd_sc_hd__o21ai_2 _6863_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_0__leaf__3035_),
    .Y(_0016_));
 sky130_fd_sc_hd__o21ai_2 _6864_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_1__leaf__3035_),
    .Y(_0017_));
 sky130_fd_sc_hd__o21ai_2 _6865_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_1__leaf__3035_),
    .Y(_0018_));
 sky130_fd_sc_hd__o21ai_2 _6866_ (.A1(_3033_),
    .A2(_3034_),
    .B1(clknet_1_1__leaf__3035_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_4 _6867_ (.A(_3024_),
    .X(_3036_));
 sky130_fd_sc_hd__buf_4 _6868_ (.A(_3027_),
    .X(_3037_));
 sky130_fd_sc_hd__buf_1 _6869_ (.A(clknet_1_0__leaf__3031_),
    .X(_3038_));
 sky130_fd_sc_hd__o21ai_2 _6870_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_1__leaf__3038_),
    .Y(_0020_));
 sky130_fd_sc_hd__o21ai_2 _6871_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_1__leaf__3038_),
    .Y(_0021_));
 sky130_fd_sc_hd__o21ai_2 _6872_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_1__leaf__3038_),
    .Y(_0022_));
 sky130_fd_sc_hd__o21ai_2 _6873_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_1__leaf__3038_),
    .Y(_0023_));
 sky130_fd_sc_hd__o21ai_2 _6874_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_0__leaf__3038_),
    .Y(_0024_));
 sky130_fd_sc_hd__o21ai_2 _6875_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_0__leaf__3038_),
    .Y(_0025_));
 sky130_fd_sc_hd__o21ai_2 _6876_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_0__leaf__3038_),
    .Y(_0026_));
 sky130_fd_sc_hd__o21ai_2 _6877_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_0__leaf__3038_),
    .Y(_0027_));
 sky130_fd_sc_hd__o21ai_2 _6878_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_0__leaf__3038_),
    .Y(_0028_));
 sky130_fd_sc_hd__o21ai_2 _6879_ (.A1(_3036_),
    .A2(_3037_),
    .B1(clknet_1_0__leaf__3038_),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_4 _6880_ (.A(_3024_),
    .X(_3039_));
 sky130_fd_sc_hd__buf_4 _6881_ (.A(_3027_),
    .X(_3040_));
 sky130_fd_sc_hd__buf_1 _6882_ (.A(clknet_1_0__leaf__3031_),
    .X(_3041_));
 sky130_fd_sc_hd__o21ai_2 _6883_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_1__leaf__3041_),
    .Y(_0030_));
 sky130_fd_sc_hd__o21ai_2 _6884_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_1__leaf__3041_),
    .Y(_0031_));
 sky130_fd_sc_hd__o21ai_2 _6885_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_1__leaf__3041_),
    .Y(_0032_));
 sky130_fd_sc_hd__o21ai_2 _6886_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_0__leaf__3041_),
    .Y(_0033_));
 sky130_fd_sc_hd__o21ai_2 _6887_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_1__leaf__3041_),
    .Y(_0034_));
 sky130_fd_sc_hd__o21ai_2 _6888_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_0__leaf__3041_),
    .Y(_0035_));
 sky130_fd_sc_hd__o21ai_2 _6889_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_1__leaf__3041_),
    .Y(_0036_));
 sky130_fd_sc_hd__o21ai_2 _6890_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_1__leaf__3041_),
    .Y(_0037_));
 sky130_fd_sc_hd__o21ai_2 _6891_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_0__leaf__3041_),
    .Y(_0038_));
 sky130_fd_sc_hd__o21ai_2 _6892_ (.A1(_3039_),
    .A2(_3040_),
    .B1(clknet_1_0__leaf__3041_),
    .Y(_0039_));
 sky130_fd_sc_hd__buf_4 _6893_ (.A(_3024_),
    .X(_3042_));
 sky130_fd_sc_hd__buf_4 _6894_ (.A(_3027_),
    .X(_3043_));
 sky130_fd_sc_hd__buf_1 _6895_ (.A(clknet_1_0__leaf__3031_),
    .X(_3044_));
 sky130_fd_sc_hd__o21ai_2 _6896_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_1__leaf__3044_),
    .Y(_0040_));
 sky130_fd_sc_hd__o21ai_2 _6897_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_1__leaf__3044_),
    .Y(_0041_));
 sky130_fd_sc_hd__o21ai_2 _6898_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_1__leaf__3044_),
    .Y(_0042_));
 sky130_fd_sc_hd__o21ai_2 _6899_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_1__leaf__3044_),
    .Y(_0043_));
 sky130_fd_sc_hd__o21ai_2 _6900_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_0__leaf__3044_),
    .Y(_0044_));
 sky130_fd_sc_hd__o21ai_2 _6901_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_0__leaf__3044_),
    .Y(_0045_));
 sky130_fd_sc_hd__o21ai_2 _6902_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_0__leaf__3044_),
    .Y(_0046_));
 sky130_fd_sc_hd__o21ai_2 _6903_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_0__leaf__3044_),
    .Y(_0047_));
 sky130_fd_sc_hd__o21ai_2 _6904_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_0__leaf__3044_),
    .Y(_0048_));
 sky130_fd_sc_hd__o21ai_2 _6905_ (.A1(_3042_),
    .A2(_3043_),
    .B1(clknet_1_0__leaf__3044_),
    .Y(_0049_));
 sky130_fd_sc_hd__buf_4 _6906_ (.A(_3024_),
    .X(_3045_));
 sky130_fd_sc_hd__buf_4 _6907_ (.A(_3027_),
    .X(_3046_));
 sky130_fd_sc_hd__buf_1 _6908_ (.A(clknet_1_1__leaf__3031_),
    .X(_3047_));
 sky130_fd_sc_hd__o21ai_2 _6909_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_0__leaf__3047_),
    .Y(_0050_));
 sky130_fd_sc_hd__o21ai_2 _6910_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_0__leaf__3047_),
    .Y(_0051_));
 sky130_fd_sc_hd__o21ai_2 _6911_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_0__leaf__3047_),
    .Y(_0052_));
 sky130_fd_sc_hd__o21ai_2 _6912_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_0__leaf__3047_),
    .Y(_0053_));
 sky130_fd_sc_hd__o21ai_2 _6913_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_1__leaf__3047_),
    .Y(_0054_));
 sky130_fd_sc_hd__o21ai_2 _6914_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_1__leaf__3047_),
    .Y(_0055_));
 sky130_fd_sc_hd__o21ai_2 _6915_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_1__leaf__3047_),
    .Y(_0056_));
 sky130_fd_sc_hd__o21ai_2 _6916_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_1__leaf__3047_),
    .Y(_0057_));
 sky130_fd_sc_hd__o21ai_2 _6917_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_1__leaf__3047_),
    .Y(_0058_));
 sky130_fd_sc_hd__o21ai_2 _6918_ (.A1(_3045_),
    .A2(_3046_),
    .B1(clknet_1_1__leaf__3047_),
    .Y(_0059_));
 sky130_fd_sc_hd__buf_4 _6919_ (.A(_3024_),
    .X(_3048_));
 sky130_fd_sc_hd__buf_4 _6920_ (.A(_3027_),
    .X(_3049_));
 sky130_fd_sc_hd__buf_1 _6921_ (.A(clknet_1_1__leaf__3031_),
    .X(_3050_));
 sky130_fd_sc_hd__o21ai_2 _6922_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_0__leaf__3050_),
    .Y(_0060_));
 sky130_fd_sc_hd__o21ai_2 _6923_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_0__leaf__3050_),
    .Y(_0061_));
 sky130_fd_sc_hd__o21ai_2 _6924_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_0__leaf__3050_),
    .Y(_0062_));
 sky130_fd_sc_hd__o21ai_2 _6925_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_0__leaf__3050_),
    .Y(_0063_));
 sky130_fd_sc_hd__o21ai_2 _6926_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_1__leaf__3050_),
    .Y(_0064_));
 sky130_fd_sc_hd__o21ai_2 _6927_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_0__leaf__3050_),
    .Y(_0065_));
 sky130_fd_sc_hd__o21ai_2 _6928_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_1__leaf__3050_),
    .Y(_0066_));
 sky130_fd_sc_hd__o21ai_2 _6929_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_1__leaf__3050_),
    .Y(_0067_));
 sky130_fd_sc_hd__o21ai_2 _6930_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_1__leaf__3050_),
    .Y(_0068_));
 sky130_fd_sc_hd__o21ai_2 _6931_ (.A1(_3048_),
    .A2(_3049_),
    .B1(clknet_1_1__leaf__3050_),
    .Y(_0069_));
 sky130_fd_sc_hd__buf_4 _6932_ (.A(_3024_),
    .X(_3051_));
 sky130_fd_sc_hd__buf_4 _6933_ (.A(_3027_),
    .X(_3052_));
 sky130_fd_sc_hd__buf_1 _6934_ (.A(clknet_1_1__leaf__3031_),
    .X(_3053_));
 sky130_fd_sc_hd__o21ai_2 _6935_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_0__leaf__3053_),
    .Y(_0070_));
 sky130_fd_sc_hd__o21ai_2 _6936_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_0__leaf__3053_),
    .Y(_0071_));
 sky130_fd_sc_hd__o21ai_2 _6937_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_0__leaf__3053_),
    .Y(_0072_));
 sky130_fd_sc_hd__o21ai_2 _6938_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_0__leaf__3053_),
    .Y(_0073_));
 sky130_fd_sc_hd__o21ai_2 _6939_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_0__leaf__3053_),
    .Y(_0074_));
 sky130_fd_sc_hd__o21ai_2 _6940_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_0__leaf__3053_),
    .Y(_0075_));
 sky130_fd_sc_hd__o21ai_2 _6941_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_1__leaf__3053_),
    .Y(_0076_));
 sky130_fd_sc_hd__o21ai_2 _6942_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_1__leaf__3053_),
    .Y(_0077_));
 sky130_fd_sc_hd__o21ai_2 _6943_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_1__leaf__3053_),
    .Y(_0078_));
 sky130_fd_sc_hd__o21ai_2 _6944_ (.A1(_3051_),
    .A2(_3052_),
    .B1(clknet_1_1__leaf__3053_),
    .Y(_0079_));
 sky130_fd_sc_hd__buf_4 _6945_ (.A(_3024_),
    .X(_3054_));
 sky130_fd_sc_hd__buf_4 _6946_ (.A(_3027_),
    .X(_3055_));
 sky130_fd_sc_hd__buf_1 _6947_ (.A(clknet_1_1__leaf__3031_),
    .X(_3056_));
 sky130_fd_sc_hd__o21ai_2 _6948_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_0__leaf__3056_),
    .Y(_0080_));
 sky130_fd_sc_hd__o21ai_2 _6949_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_0__leaf__3056_),
    .Y(_0081_));
 sky130_fd_sc_hd__o21ai_2 _6950_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_0__leaf__3056_),
    .Y(_0082_));
 sky130_fd_sc_hd__o21ai_2 _6951_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_0__leaf__3056_),
    .Y(_0083_));
 sky130_fd_sc_hd__o21ai_2 _6952_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_1__leaf__3056_),
    .Y(_0084_));
 sky130_fd_sc_hd__o21ai_2 _6953_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_1__leaf__3056_),
    .Y(_0085_));
 sky130_fd_sc_hd__o21ai_2 _6954_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_1__leaf__3056_),
    .Y(_0086_));
 sky130_fd_sc_hd__o21ai_2 _6955_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_1__leaf__3056_),
    .Y(_0087_));
 sky130_fd_sc_hd__o21ai_2 _6956_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_1__leaf__3056_),
    .Y(_0088_));
 sky130_fd_sc_hd__o21ai_2 _6957_ (.A1(_3054_),
    .A2(_3055_),
    .B1(clknet_1_1__leaf__3056_),
    .Y(_0089_));
 sky130_fd_sc_hd__buf_4 _6958_ (.A(_3023_),
    .X(_3057_));
 sky130_fd_sc_hd__buf_4 _6959_ (.A(_3026_),
    .X(_3058_));
 sky130_fd_sc_hd__buf_1 _6960_ (.A(clknet_1_1__leaf__3030_),
    .X(_3059_));
 sky130_fd_sc_hd__o21ai_2 _6961_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_1__leaf__3059_),
    .Y(_0090_));
 sky130_fd_sc_hd__o21ai_2 _6962_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_0__leaf__3059_),
    .Y(_0091_));
 sky130_fd_sc_hd__o21ai_2 _6963_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_1__leaf__3059_),
    .Y(_0092_));
 sky130_fd_sc_hd__o21ai_2 _6964_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_1__leaf__3059_),
    .Y(_0093_));
 sky130_fd_sc_hd__o21ai_2 _6965_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_0__leaf__3059_),
    .Y(_0094_));
 sky130_fd_sc_hd__o21ai_2 _6966_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_1__leaf__3059_),
    .Y(_0095_));
 sky130_fd_sc_hd__o21ai_2 _6967_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_1__leaf__3059_),
    .Y(_0096_));
 sky130_fd_sc_hd__o21ai_2 _6968_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_0__leaf__3059_),
    .Y(_0097_));
 sky130_fd_sc_hd__o21ai_2 _6969_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_0__leaf__3059_),
    .Y(_0098_));
 sky130_fd_sc_hd__o21ai_2 _6970_ (.A1(_3057_),
    .A2(_3058_),
    .B1(clknet_1_0__leaf__3059_),
    .Y(_0099_));
 sky130_fd_sc_hd__buf_4 _6971_ (.A(_3023_),
    .X(_3060_));
 sky130_fd_sc_hd__buf_4 _6972_ (.A(_3026_),
    .X(_3061_));
 sky130_fd_sc_hd__buf_1 _6973_ (.A(clknet_1_1__leaf__3030_),
    .X(_3062_));
 sky130_fd_sc_hd__o21ai_2 _6974_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_1__leaf__3062_),
    .Y(_0100_));
 sky130_fd_sc_hd__o21ai_2 _6975_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_1__leaf__3062_),
    .Y(_0101_));
 sky130_fd_sc_hd__o21ai_2 _6976_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_1__leaf__3062_),
    .Y(_0102_));
 sky130_fd_sc_hd__o21ai_2 _6977_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_1__leaf__3062_),
    .Y(_0103_));
 sky130_fd_sc_hd__o21ai_2 _6978_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_0__leaf__3062_),
    .Y(_0104_));
 sky130_fd_sc_hd__o21ai_2 _6979_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_1__leaf__3062_),
    .Y(_0105_));
 sky130_fd_sc_hd__o21ai_2 _6980_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_0__leaf__3062_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ai_2 _6981_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_0__leaf__3062_),
    .Y(_0107_));
 sky130_fd_sc_hd__o21ai_2 _6982_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_0__leaf__3062_),
    .Y(_0108_));
 sky130_fd_sc_hd__o21ai_2 _6983_ (.A1(_3060_),
    .A2(_3061_),
    .B1(clknet_1_0__leaf__3062_),
    .Y(_0109_));
 sky130_fd_sc_hd__buf_4 _6984_ (.A(_3023_),
    .X(_3063_));
 sky130_fd_sc_hd__buf_4 _6985_ (.A(_3026_),
    .X(_3064_));
 sky130_fd_sc_hd__buf_1 _6986_ (.A(clknet_1_1__leaf__3030_),
    .X(_3065_));
 sky130_fd_sc_hd__o21ai_2 _6987_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_0__leaf__3065_),
    .Y(_0110_));
 sky130_fd_sc_hd__o21ai_2 _6988_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_0__leaf__3065_),
    .Y(_0111_));
 sky130_fd_sc_hd__o21ai_2 _6989_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_1__leaf__3065_),
    .Y(_0112_));
 sky130_fd_sc_hd__o21ai_2 _6990_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_1__leaf__3065_),
    .Y(_0113_));
 sky130_fd_sc_hd__o21ai_2 _6991_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_1__leaf__3065_),
    .Y(_0114_));
 sky130_fd_sc_hd__o21ai_2 _6992_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_0__leaf__3065_),
    .Y(_0115_));
 sky130_fd_sc_hd__o21ai_2 _6993_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_1__leaf__3065_),
    .Y(_0116_));
 sky130_fd_sc_hd__o21ai_2 _6994_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_1__leaf__3065_),
    .Y(_0117_));
 sky130_fd_sc_hd__o21ai_2 _6995_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_1__leaf__3065_),
    .Y(_0118_));
 sky130_fd_sc_hd__o21ai_2 _6996_ (.A1(_3063_),
    .A2(_3064_),
    .B1(clknet_1_0__leaf__3065_),
    .Y(_0119_));
 sky130_fd_sc_hd__buf_4 _6997_ (.A(_3023_),
    .X(_3066_));
 sky130_fd_sc_hd__buf_4 _6998_ (.A(_3026_),
    .X(_3067_));
 sky130_fd_sc_hd__buf_1 _6999_ (.A(clknet_1_0__leaf__3030_),
    .X(_3068_));
 sky130_fd_sc_hd__o21ai_2 _7000_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_1__leaf__3068_),
    .Y(_0120_));
 sky130_fd_sc_hd__o21ai_2 _7001_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_1__leaf__3068_),
    .Y(_0121_));
 sky130_fd_sc_hd__o21ai_2 _7002_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_0__leaf__3068_),
    .Y(_0122_));
 sky130_fd_sc_hd__o21ai_2 _7003_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_0__leaf__3068_),
    .Y(_0123_));
 sky130_fd_sc_hd__o21ai_2 _7004_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_1__leaf__3068_),
    .Y(_0124_));
 sky130_fd_sc_hd__o21ai_2 _7005_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_0__leaf__3068_),
    .Y(_0125_));
 sky130_fd_sc_hd__o21ai_2 _7006_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_0__leaf__3068_),
    .Y(_0126_));
 sky130_fd_sc_hd__o21ai_2 _7007_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_0__leaf__3068_),
    .Y(_0127_));
 sky130_fd_sc_hd__o21ai_2 _7008_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_1__leaf__3068_),
    .Y(_0128_));
 sky130_fd_sc_hd__o21ai_2 _7009_ (.A1(_3066_),
    .A2(_3067_),
    .B1(clknet_1_1__leaf__3068_),
    .Y(_0129_));
 sky130_fd_sc_hd__clkbuf_8 _7010_ (.A(_3023_),
    .X(_3069_));
 sky130_fd_sc_hd__buf_4 _7011_ (.A(_3026_),
    .X(_3070_));
 sky130_fd_sc_hd__buf_1 _7012_ (.A(clknet_1_0__leaf__3030_),
    .X(_3071_));
 sky130_fd_sc_hd__o21ai_2 _7013_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_1__leaf__3071_),
    .Y(_0130_));
 sky130_fd_sc_hd__o21ai_2 _7014_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_0__leaf__3071_),
    .Y(_0131_));
 sky130_fd_sc_hd__o21ai_2 _7015_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_0__leaf__3071_),
    .Y(_0132_));
 sky130_fd_sc_hd__o21ai_2 _7016_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_0__leaf__3071_),
    .Y(_0133_));
 sky130_fd_sc_hd__o21ai_2 _7017_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_0__leaf__3071_),
    .Y(_0134_));
 sky130_fd_sc_hd__o21ai_2 _7018_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_0__leaf__3071_),
    .Y(_0135_));
 sky130_fd_sc_hd__o21ai_2 _7019_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_0__leaf__3071_),
    .Y(_0136_));
 sky130_fd_sc_hd__o21ai_2 _7020_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_1__leaf__3071_),
    .Y(_0137_));
 sky130_fd_sc_hd__o21ai_2 _7021_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_1__leaf__3071_),
    .Y(_0138_));
 sky130_fd_sc_hd__o21ai_2 _7022_ (.A1(_3069_),
    .A2(_3070_),
    .B1(clknet_1_1__leaf__3071_),
    .Y(_0139_));
 sky130_fd_sc_hd__buf_4 _7023_ (.A(_3023_),
    .X(_3072_));
 sky130_fd_sc_hd__buf_4 _7024_ (.A(_3026_),
    .X(_3073_));
 sky130_fd_sc_hd__buf_1 _7025_ (.A(clknet_1_0__leaf__3030_),
    .X(_3074_));
 sky130_fd_sc_hd__o21ai_2 _7026_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_1__leaf__3074_),
    .Y(_0140_));
 sky130_fd_sc_hd__o21ai_2 _7027_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_1__leaf__3074_),
    .Y(_0141_));
 sky130_fd_sc_hd__o21ai_2 _7028_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_0__leaf__3074_),
    .Y(_0142_));
 sky130_fd_sc_hd__o21ai_2 _7029_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_1__leaf__3074_),
    .Y(_0143_));
 sky130_fd_sc_hd__o21ai_2 _7030_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_1__leaf__3074_),
    .Y(_0144_));
 sky130_fd_sc_hd__o21ai_2 _7031_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_0__leaf__3074_),
    .Y(_0145_));
 sky130_fd_sc_hd__o21ai_2 _7032_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_0__leaf__3074_),
    .Y(_0146_));
 sky130_fd_sc_hd__o21ai_2 _7033_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_0__leaf__3074_),
    .Y(_0147_));
 sky130_fd_sc_hd__o21ai_2 _7034_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_0__leaf__3074_),
    .Y(_0148_));
 sky130_fd_sc_hd__o21ai_2 _7035_ (.A1(_3072_),
    .A2(_3073_),
    .B1(clknet_1_0__leaf__3074_),
    .Y(_0149_));
 sky130_fd_sc_hd__buf_4 _7036_ (.A(_3023_),
    .X(_3075_));
 sky130_fd_sc_hd__buf_4 _7037_ (.A(_3026_),
    .X(_3076_));
 sky130_fd_sc_hd__buf_1 _7038_ (.A(clknet_1_0__leaf__3030_),
    .X(_3077_));
 sky130_fd_sc_hd__o21ai_2 _7039_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_1__leaf__3077_),
    .Y(_0150_));
 sky130_fd_sc_hd__o21ai_2 _7040_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_1__leaf__3077_),
    .Y(_0151_));
 sky130_fd_sc_hd__o21ai_2 _7041_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_1__leaf__3077_),
    .Y(_0152_));
 sky130_fd_sc_hd__o21ai_2 _7042_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_1__leaf__3077_),
    .Y(_0153_));
 sky130_fd_sc_hd__o21ai_2 _7043_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_0__leaf__3077_),
    .Y(_0154_));
 sky130_fd_sc_hd__o21ai_2 _7044_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_0__leaf__3077_),
    .Y(_0155_));
 sky130_fd_sc_hd__o21ai_2 _7045_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_0__leaf__3077_),
    .Y(_0156_));
 sky130_fd_sc_hd__o21ai_2 _7046_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_0__leaf__3077_),
    .Y(_0157_));
 sky130_fd_sc_hd__o21ai_2 _7047_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_0__leaf__3077_),
    .Y(_0158_));
 sky130_fd_sc_hd__o21ai_2 _7048_ (.A1(_3075_),
    .A2(_3076_),
    .B1(clknet_1_0__leaf__3077_),
    .Y(_0159_));
 sky130_fd_sc_hd__o21ai_2 _7049_ (.A1(_3024_),
    .A2(_3027_),
    .B1(clknet_1_0__leaf__3031_),
    .Y(_0160_));
 sky130_fd_sc_hd__dfxtp_1 _7050_ (.CLK(_0000_),
    .D(_0161_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfxtp_1 _7051_ (.CLK(_0001_),
    .D(_0162_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfxtp_1 _7052_ (.CLK(_0002_),
    .D(_0163_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfxtp_1 _7053_ (.CLK(_0003_),
    .D(_0164_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfxtp_1 _7054_ (.CLK(_0004_),
    .D(_0165_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfxtp_1 _7055_ (.CLK(_0005_),
    .D(_0166_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfxtp_1 _7056_ (.CLK(_0006_),
    .D(_0167_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfxtp_1 _7057_ (.CLK(_0007_),
    .D(_0168_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfxtp_1 _7058_ (.CLK(_0008_),
    .D(_0169_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfxtp_1 _7059_ (.CLK(_0009_),
    .D(_0170_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfxtp_1 _7060_ (.CLK(_0010_),
    .D(_0171_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfxtp_2 _7061_ (.CLK(_0011_),
    .D(_0172_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfxtp_1 _7062_ (.CLK(_0012_),
    .D(_0173_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfxtp_1 _7063_ (.CLK(_0013_),
    .D(_0174_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfxtp_1 _7064_ (.CLK(_0014_),
    .D(_0175_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfxtp_2 _7065_ (.CLK(_0015_),
    .D(_0176_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_1 _7066_ (.CLK(_0016_),
    .D(_0177_),
    .Q(\egd_top.BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7067_ (.CLK(_0017_),
    .D(_0178_),
    .Q(\egd_top.BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7068_ (.CLK(_0018_),
    .D(_0179_),
    .Q(\egd_top.BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7069_ (.CLK(_0019_),
    .D(_0180_),
    .Q(\egd_top.BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7070_ (.CLK(_0020_),
    .D(_0181_),
    .Q(\egd_top.BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7071_ (.CLK(_0021_),
    .D(_0182_),
    .Q(\egd_top.BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7072_ (.CLK(_0022_),
    .D(_0183_),
    .Q(\egd_top.BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7073_ (.CLK(_0023_),
    .D(_0184_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfxtp_1 _7074_ (.CLK(_0024_),
    .D(_0185_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfxtp_1 _7075_ (.CLK(_0025_),
    .D(_0186_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfxtp_2 _7076_ (.CLK(_0026_),
    .D(_0187_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfxtp_1 _7077_ (.CLK(_0027_),
    .D(_0188_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfxtp_1 _7078_ (.CLK(_0028_),
    .D(_0189_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfxtp_1 _7079_ (.CLK(_0029_),
    .D(_0190_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfxtp_1 _7080_ (.CLK(_0030_),
    .D(_0191_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfxtp_1 _7081_ (.CLK(_0031_),
    .D(_0192_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfxtp_1 _7082_ (.CLK(_0032_),
    .D(_0193_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfxtp_1 _7083_ (.CLK(_0033_),
    .D(_0194_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfxtp_1 _7084_ (.CLK(_0034_),
    .D(_0195_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfxtp_1 _7085_ (.CLK(_0035_),
    .D(_0196_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfxtp_1 _7086_ (.CLK(_0036_),
    .D(_0197_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfxtp_1 _7087_ (.CLK(_0037_),
    .D(_0198_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfxtp_1 _7088_ (.CLK(_0038_),
    .D(_0199_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfxtp_1 _7089_ (.CLK(_0039_),
    .D(_0200_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfxtp_1 _7090_ (.CLK(_0040_),
    .D(_0201_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfxtp_1 _7091_ (.CLK(_0041_),
    .D(_0202_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfxtp_1 _7092_ (.CLK(_0042_),
    .D(_0203_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfxtp_1 _7093_ (.CLK(_0043_),
    .D(_0204_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfxtp_1 _7094_ (.CLK(_0044_),
    .D(_0205_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfxtp_1 _7095_ (.CLK(_0045_),
    .D(_0206_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _7096_ (.CLK(_0046_),
    .D(_0207_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_2 _7097_ (.CLK(_0047_),
    .D(_0208_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _7098_ (.CLK(_0048_),
    .D(_0209_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _7099_ (.CLK(_0049_),
    .D(_0210_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _7100_ (.CLK(_0050_),
    .D(_0211_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _7101_ (.CLK(_0051_),
    .D(_0212_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _7102_ (.CLK(_0052_),
    .D(_0213_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _7103_ (.CLK(_0053_),
    .D(_0214_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _7104_ (.CLK(_0054_),
    .D(_0215_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _7105_ (.CLK(_0055_),
    .D(_0216_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _7106_ (.CLK(_0056_),
    .D(_0217_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _7107_ (.CLK(_0057_),
    .D(_0218_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _7108_ (.CLK(_0058_),
    .D(_0219_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _7109_ (.CLK(_0059_),
    .D(_0220_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _7110_ (.CLK(_0060_),
    .D(_0221_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _7111_ (.CLK(_0061_),
    .D(_0222_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _7112_ (.CLK(_0062_),
    .D(_0223_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _7113_ (.CLK(_0063_),
    .D(_0224_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_2 _7114_ (.CLK(_0064_),
    .D(_0225_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _7115_ (.CLK(_0065_),
    .D(_0226_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _7116_ (.CLK(_0066_),
    .D(_0227_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _7117_ (.CLK(_0067_),
    .D(_0228_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _7118_ (.CLK(_0068_),
    .D(_0229_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _7119_ (.CLK(_0069_),
    .D(_0230_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _7120_ (.CLK(_0070_),
    .D(_0231_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _7121_ (.CLK(_0071_),
    .D(_0232_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _7122_ (.CLK(_0072_),
    .D(_0233_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _7123_ (.CLK(_0073_),
    .D(_0234_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _7124_ (.CLK(_0074_),
    .D(_0235_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _7125_ (.CLK(_0075_),
    .D(_0236_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _7126_ (.CLK(_0076_),
    .D(_0237_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _7127_ (.CLK(_0077_),
    .D(_0238_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _7128_ (.CLK(_0078_),
    .D(_0239_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _7129_ (.CLK(_0079_),
    .D(_0240_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _7130_ (.CLK(_0080_),
    .D(_0241_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _7131_ (.CLK(_0081_),
    .D(_0242_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _7132_ (.CLK(_0082_),
    .D(_0243_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _7133_ (.CLK(_0083_),
    .D(_0244_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _7134_ (.CLK(_0084_),
    .D(_0245_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_2 _7135_ (.CLK(_0085_),
    .D(_0246_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _7136_ (.CLK(_0086_),
    .D(_0247_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _7137_ (.CLK(_0087_),
    .D(_0248_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _7138_ (.CLK(_0088_),
    .D(_0249_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_2 _7139_ (.CLK(_0089_),
    .D(_0250_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _7140_ (.CLK(_0090_),
    .D(_0251_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _7141_ (.CLK(_0091_),
    .D(_0252_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _7142_ (.CLK(_0092_),
    .D(_0253_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _7143_ (.CLK(_0093_),
    .D(_0254_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _7144_ (.CLK(_0094_),
    .D(_0255_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _7145_ (.CLK(_0095_),
    .D(_0256_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _7146_ (.CLK(_0096_),
    .D(_0257_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _7147_ (.CLK(_0097_),
    .D(_0258_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _7148_ (.CLK(_0098_),
    .D(_0259_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _7149_ (.CLK(_0099_),
    .D(_0260_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _7150_ (.CLK(_0100_),
    .D(_0261_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _7151_ (.CLK(_0101_),
    .D(_0262_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _7152_ (.CLK(_0102_),
    .D(_0263_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _7153_ (.CLK(_0103_),
    .D(_0264_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7154_ (.CLK(_0104_),
    .D(_0265_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7155_ (.CLK(_0105_),
    .D(_0266_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7156_ (.CLK(_0106_),
    .D(_0267_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7157_ (.CLK(_0107_),
    .D(_0268_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7158_ (.CLK(_0108_),
    .D(_0269_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7159_ (.CLK(_0109_),
    .D(_0270_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7160_ (.CLK(_0110_),
    .D(_0271_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7161_ (.CLK(_0111_),
    .D(_0272_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7162_ (.CLK(_0112_),
    .D(_0273_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7163_ (.CLK(_0113_),
    .D(_0274_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7164_ (.CLK(_0114_),
    .D(_0275_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7165_ (.CLK(_0115_),
    .D(_0276_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7166_ (.CLK(_0116_),
    .D(_0277_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7167_ (.CLK(_0117_),
    .D(_0278_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7168_ (.CLK(_0118_),
    .D(_0279_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7169_ (.CLK(_0119_),
    .D(_0280_),
    .Q(\egd_top.BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7170_ (.CLK(_0120_),
    .D(_0281_),
    .Q(\egd_top.BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7171_ (.CLK(_0121_),
    .D(_0282_),
    .Q(\egd_top.BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7172_ (.CLK(_0122_),
    .D(_0283_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7173_ (.CLK(_0123_),
    .D(_0284_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7174_ (.CLK(_0124_),
    .D(_0285_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7175_ (.CLK(_0125_),
    .D(_0286_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7176_ (.CLK(_0126_),
    .D(_0287_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7177_ (.CLK(_0127_),
    .D(_0288_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7178_ (.CLK(_0128_),
    .D(_0289_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7179_ (.CLK(_0129_),
    .D(_0290_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfxtp_2 _7180_ (.CLK(_0130_),
    .D(_0291_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7181_ (.CLK(_0131_),
    .D(_0292_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfxtp_2 _7182_ (.CLK(_0132_),
    .D(_0293_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfxtp_2 _7183_ (.CLK(_0133_),
    .D(_0294_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfxtp_2 _7184_ (.CLK(_0134_),
    .D(_0295_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7185_ (.CLK(_0135_),
    .D(_0296_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7186_ (.CLK(_0136_),
    .D(_0297_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7187_ (.CLK(_0137_),
    .D(_0298_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfxtp_1 _7188_ (.CLK(_0138_),
    .D(_0299_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfxtp_1 _7189_ (.CLK(_0139_),
    .D(_0300_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfxtp_1 _7190_ (.CLK(_0140_),
    .D(_0301_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfxtp_1 _7191_ (.CLK(_0141_),
    .D(_0302_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfxtp_1 _7192_ (.CLK(_0142_),
    .D(_0303_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfxtp_1 _7193_ (.CLK(_0143_),
    .D(_0304_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfxtp_1 _7194_ (.CLK(_0144_),
    .D(_0305_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfxtp_1 _7195_ (.CLK(_0145_),
    .D(_0306_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfxtp_1 _7196_ (.CLK(_0146_),
    .D(_0307_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfxtp_1 _7197_ (.CLK(_0147_),
    .D(_0308_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfxtp_1 _7198_ (.CLK(_0148_),
    .D(_0309_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfxtp_1 _7199_ (.CLK(_0149_),
    .D(_0310_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfxtp_1 _7200_ (.CLK(_0150_),
    .D(_0311_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfxtp_1 _7201_ (.CLK(_0151_),
    .D(_0312_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfxtp_1 _7202_ (.CLK(_0152_),
    .D(_0313_),
    .Q(\egd_top.BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfxtp_1 _7203_ (.CLK(_0153_),
    .D(_0314_),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfxtp_2 _7204_ (.CLK(_0154_),
    .D(_0315_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _7205_ (.CLK(_0155_),
    .D(_0316_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _7206_ (.CLK(_0156_),
    .D(_0317_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _7207_ (.CLK(_0157_),
    .D(_0318_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_2 _7208_ (.CLK(_0158_),
    .D(_0319_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_2 _7209_ (.CLK(_0159_),
    .D(_0320_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_2 _7210_ (.CLK(_0160_),
    .D(_0321_),
    .Q(net38));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3030_ (.A(_3030_),
    .X(clknet_0__3030_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3031_ (.A(_3031_),
    .X(clknet_0__3031_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3032_ (.A(_3032_),
    .X(clknet_0__3032_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3035_ (.A(_3035_),
    .X(clknet_0__3035_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3038_ (.A(_3038_),
    .X(clknet_0__3038_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3041_ (.A(_3041_),
    .X(clknet_0__3041_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3044_ (.A(_3044_),
    .X(clknet_0__3044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3047_ (.A(_3047_),
    .X(clknet_0__3047_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3050_ (.A(_3050_),
    .X(clknet_0__3050_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3053_ (.A(_3053_),
    .X(clknet_0__3053_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3056_ (.A(_3056_),
    .X(clknet_0__3056_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3059_ (.A(_3059_),
    .X(clknet_0__3059_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3062_ (.A(_3062_),
    .X(clknet_0__3062_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3065_ (.A(_3065_),
    .X(clknet_0__3065_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3068_ (.A(_3068_),
    .X(clknet_0__3068_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3071_ (.A(_3071_),
    .X(clknet_0__3071_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3074_ (.A(_3074_),
    .X(clknet_0__3074_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__3077_ (.A(_3077_),
    .X(clknet_0__3077_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3030_ (.A(clknet_0__3030_),
    .X(clknet_1_0__leaf__3030_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3031_ (.A(clknet_0__3031_),
    .X(clknet_1_0__leaf__3031_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3032_ (.A(clknet_0__3032_),
    .X(clknet_1_0__leaf__3032_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3035_ (.A(clknet_0__3035_),
    .X(clknet_1_0__leaf__3035_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3038_ (.A(clknet_0__3038_),
    .X(clknet_1_0__leaf__3038_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3041_ (.A(clknet_0__3041_),
    .X(clknet_1_0__leaf__3041_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3044_ (.A(clknet_0__3044_),
    .X(clknet_1_0__leaf__3044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3047_ (.A(clknet_0__3047_),
    .X(clknet_1_0__leaf__3047_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3050_ (.A(clknet_0__3050_),
    .X(clknet_1_0__leaf__3050_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3053_ (.A(clknet_0__3053_),
    .X(clknet_1_0__leaf__3053_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3056_ (.A(clknet_0__3056_),
    .X(clknet_1_0__leaf__3056_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3059_ (.A(clknet_0__3059_),
    .X(clknet_1_0__leaf__3059_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3062_ (.A(clknet_0__3062_),
    .X(clknet_1_0__leaf__3062_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3065_ (.A(clknet_0__3065_),
    .X(clknet_1_0__leaf__3065_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3068_ (.A(clknet_0__3068_),
    .X(clknet_1_0__leaf__3068_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3071_ (.A(clknet_0__3071_),
    .X(clknet_1_0__leaf__3071_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3074_ (.A(clknet_0__3074_),
    .X(clknet_1_0__leaf__3074_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__3077_ (.A(clknet_0__3077_),
    .X(clknet_1_0__leaf__3077_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3030_ (.A(clknet_0__3030_),
    .X(clknet_1_1__leaf__3030_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3031_ (.A(clknet_0__3031_),
    .X(clknet_1_1__leaf__3031_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3032_ (.A(clknet_0__3032_),
    .X(clknet_1_1__leaf__3032_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3035_ (.A(clknet_0__3035_),
    .X(clknet_1_1__leaf__3035_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3038_ (.A(clknet_0__3038_),
    .X(clknet_1_1__leaf__3038_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3041_ (.A(clknet_0__3041_),
    .X(clknet_1_1__leaf__3041_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3044_ (.A(clknet_0__3044_),
    .X(clknet_1_1__leaf__3044_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3047_ (.A(clknet_0__3047_),
    .X(clknet_1_1__leaf__3047_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3050_ (.A(clknet_0__3050_),
    .X(clknet_1_1__leaf__3050_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3053_ (.A(clknet_0__3053_),
    .X(clknet_1_1__leaf__3053_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3056_ (.A(clknet_0__3056_),
    .X(clknet_1_1__leaf__3056_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3059_ (.A(clknet_0__3059_),
    .X(clknet_1_1__leaf__3059_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3062_ (.A(clknet_0__3062_),
    .X(clknet_1_1__leaf__3062_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3065_ (.A(clknet_0__3065_),
    .X(clknet_1_1__leaf__3065_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3068_ (.A(clknet_0__3068_),
    .X(clknet_1_1__leaf__3068_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3071_ (.A(clknet_0__3071_),
    .X(clknet_1_1__leaf__3071_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3074_ (.A(clknet_0__3074_),
    .X(clknet_1_1__leaf__3074_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__3077_ (.A(clknet_0__3077_),
    .X(clknet_1_1__leaf__3077_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 hold4 (.A(net48),
    .X(net42));
 sky130_fd_sc_hd__buf_2 hold5 (.A(_2655_),
    .X(net43));
 sky130_fd_sc_hd__buf_1 hold6 (.A(\egd_top.BitStream_buffer.buffer_index[5] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_3125_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input1 (.A(la_data_in_47_32[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(la_data_in_47_32[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(la_data_in_47_32[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(la_data_in_47_32[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(la_data_in_47_32[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(la_data_in_47_32[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(la_data_in_47_32[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(la_data_in_47_32[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(la_data_in_49_48[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(la_data_in_49_48[1]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(la_data_in_64),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(la_data_in_47_32[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(la_data_in_65),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(la_oenb_64),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(la_oenb_65),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input23 (.A(wb_rst_i),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input3 (.A(la_data_in_47_32[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(la_data_in_47_32[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(la_data_in_47_32[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(la_data_in_47_32[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(la_data_in_47_32[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(la_data_in_47_32[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(la_data_in_47_32[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(la_data_out_15_8[0]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(la_data_out_15_8[1]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(la_data_out_15_8[2]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_data_out_15_8[3]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(la_data_out_15_8[4]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(la_data_out_15_8[5]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(la_data_out_15_8[6]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(la_data_out_15_8[7]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(la_data_out_18_16[0]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(la_data_out_18_16[1]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(la_data_out_18_16[2]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(la_data_out_22_19[0]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(la_data_out_22_19[1]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(la_data_out_22_19[2]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(la_data_out_22_19[3]));
 sky130_fd_sc_hd__buf_2 split1 (.A(_3165_),
    .X(net39));
endmodule

