* NGSPICE file created from egd_top_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

.subckt egd_top_wrapper la_data_in_47_32[0] la_data_in_47_32[10] la_data_in_47_32[11]
+ la_data_in_47_32[12] la_data_in_47_32[13] la_data_in_47_32[14] la_data_in_47_32[15]
+ la_data_in_47_32[1] la_data_in_47_32[2] la_data_in_47_32[3] la_data_in_47_32[4]
+ la_data_in_47_32[5] la_data_in_47_32[6] la_data_in_47_32[7] la_data_in_47_32[8]
+ la_data_in_47_32[9] la_data_in_49_48[0] la_data_in_49_48[1] la_data_in_64 la_data_in_65
+ la_data_out_15_8[0] la_data_out_15_8[1] la_data_out_15_8[2] la_data_out_15_8[3]
+ la_data_out_15_8[4] la_data_out_15_8[5] la_data_out_15_8[6] la_data_out_15_8[7]
+ la_data_out_18_16[0] la_data_out_18_16[1] la_data_out_18_16[2] la_data_out_22_19[0]
+ la_data_out_22_19[1] la_data_out_22_19[2] la_data_out_22_19[3] la_oenb_64 la_oenb_65
+ vccd1 vssd1 wb_clk_i wb_rst_i
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6914_ _3045_ _3046_ clknet_1_1__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6845_ _3025_ _3028_ clknet_1_1__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3988_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__clkbuf_2
X_6776_ _2879_ _2906_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__nor2_1
X_5727_ _0877_ _0426_ _2057_ _2058_ _2059_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_60_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5658_ _0836_ _3253_ _3449_ _3257_ _1990_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__a221oi_1
X_4609_ _0800_ _0950_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__nor2_1
X_5589_ _1291_ _0366_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4960_ _3497_ _0376_ _0701_ _0379_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4891_ _3245_ _0801_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__nand2_1
X_3911_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _3449_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6630_ _2809_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__inv_2
X_3842_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _3380_ sky130_fd_sc_hd__buf_2
X_6561_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1 vccd1 vccd1
+ _2762_ sky130_fd_sc_hd__inv_2
X_3773_ egd_top.BitStream_buffer.BS_buffer\[24\] vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__inv_2
X_5512_ _1845_ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6492_ _2708_ _2689_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5443_ _1776_ _1777_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__nand2_1
X_5374_ _0509_ _0534_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nand2_1
X_7113_ _0063_ _0224_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
X_4325_ _0666_ _3368_ _0667_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7044_ _3075_ _3076_ clknet_1_0__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__o21ai_2
X_4256_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__buf_2
X_4187_ _0530_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6828_ _3017_ _3018_ vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6759_ _2946_ _2801_ _2947_ _2951_ _2952_ vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__o32a_1
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4110_ _3289_ _0406_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__and2_1
X_5090_ _0701_ _0376_ _0695_ _0379_ _1427_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4041_ _0384_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__buf_2
X_5992_ _0437_ _0527_ _0743_ _0530_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__o22ai_1
X_4943_ _3508_ _3296_ _3511_ _3246_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4874_ _1073_ _0576_ _1210_ _0580_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__a221oi_1
X_6613_ _2810_ _2760_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3825_ _3292_ _3323_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__and2_1
X_3756_ _3293_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__clkbuf_2
X_6544_ _2743_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6475_ _3218_ _3090_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3687_ _3117_ egd_top.BitStream_buffer.pc\[2\] _3216_ vssd1 vssd1 vccd1 vccd1 _3225_
+ sky130_fd_sc_hd__and3_1
X_5426_ _3380_ _3361_ _3322_ _3365_ _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a221oi_1
X_5357_ _0404_ _0427_ _1690_ _1691_ _1692_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__o2111a_1
X_4308_ _0649_ _3291_ _0650_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__o21ai_1
X_5288_ _0653_ _3291_ _1623_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__o21ai_1
X_4239_ _0582_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__buf_2
X_7027_ _3072_ _3073_ clknet_1_1__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4590_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__clkbuf_4
X_3610_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__clkbuf_4
X_3541_ _3094_ _3099_ _3089_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ _2553_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6191_ _2505_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__clkbuf_1
X_5211_ _0380_ _0351_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__nor2_1
X_5142_ _0781_ _0614_ _0932_ _0618_ _1479_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__a221oi_1
X_5073_ _3288_ _3502_ _0649_ _3505_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__o22ai_1
X_4024_ _3283_ _0344_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5975_ _2304_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4926_ _1115_ _3424_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4857_ _0509_ _0518_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3808_ _3345_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__clkbuf_2
X_6527_ net10 _0768_ _2706_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__mux2_1
X_4788_ _0976_ _3424_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__o21ai_1
X_3739_ _3276_ _3216_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__nand2_4
X_6458_ _3079_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__buf_2
X_5409_ _3270_ _1130_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__nand2_1
X_6389_ _2641_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5760_ _0605_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _2093_
+ sky130_fd_sc_hd__nand2_1
X_4711_ _1032_ _1051_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__nand2_1
X_5691_ _2013_ _2016_ _2019_ _2023_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4642_ _3327_ _3379_ _3336_ _3383_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _0509_ _0765_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3524_ _3081_ _3085_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6312_ _2588_ _2580_ vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__and2_1
X_6243_ _2541_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
X_6174_ net16 _3476_ _2480_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__mux2_1
X_5125_ _1334_ _0544_ _1462_ _0547_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5056_ _3427_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _1394_
+ sky130_fd_sc_hd__nand2_1
X_4007_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5958_ _3208_ _0360_ _0634_ _0363_ _2288_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__a221oi_1
X_4909_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5889_ _2206_ _2220_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_5 _3467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__3032_ clknet_0__3032_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3032_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6930_ _3048_ _3049_ clknet_1_1__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6861_ _3033_ _3034_ clknet_1_1__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6792_ _2983_ _2984_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__nand2_1
X_5812_ _2142_ _2143_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__nand2_1
X_5743_ _0522_ _0493_ _0495_ _0768_ _2075_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5674_ _3385_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _2007_
+ sky130_fd_sc_hd__nand2_1
X_4625_ _3264_ _3305_ _3250_ _3310_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4556_ _0451_ _0739_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4487_ _0827_ _3368_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__o21ai_1
X_6226_ _2513_ _2529_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__and2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _2482_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _0475_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _1446_
+ sky130_fd_sc_hd__nand2_1
X_6088_ _0416_ _3199_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__nand2_1
X_5039_ _0593_ _3326_ _0597_ _3330_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[7] sky130_fd_sc_hd__buf_12
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4410_ _0751_ _0752_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__nand2_1
X_5390_ _0606_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _1726_
+ sky130_fd_sc_hd__nand2_1
X_4341_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7060_ _0010_ _0171_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_4272_ _3307_ _0553_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__and2_1
X_6011_ _2327_ _2341_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__nand2_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6913_ _3045_ _3046_ clknet_1_1__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6844_ _3025_ _3028_ clknet_1_1__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3987_ _3302_ _3469_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6775_ _2965_ _2967_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5726_ _0365_ _0438_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5657_ _1988_ _1989_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__nand2_1
X_4608_ _3212_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nor2_1
X_5588_ _0369_ _3195_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4539_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6209_ _2518_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
X_7189_ _0139_ _0300_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4890_ _3237_ _3300_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__nand2_1
X_3910_ _3432_ _3435_ _3438_ _3439_ _3447_ vssd1 vssd1 vccd1 vccd1 _3448_ sky130_fd_sc_hd__a221oi_1
X_3841_ _3378_ vssd1 vssd1 vccd1 vccd1 _3379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3772_ _3309_ vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__buf_2
X_6560_ _2759_ _2760_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__nand2_1
X_5511_ _0588_ _1192_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6491_ net7 _0781_ _2707_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__mux2_1
X_5442_ _3463_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _1777_
+ sky130_fd_sc_hd__nand2_1
X_5373_ egd_top.BitStream_buffer.BS_buffer\[88\] _0494_ _0496_ _0916_ _1708_ vssd1
+ vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__a221oi_1
X_7112_ _0062_ _0223_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_4324_ _3371_ _3358_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__nand2_1
X_7043_ _3075_ _3076_ clknet_1_0__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__o21ai_2
X_4255_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__clkbuf_2
X_4186_ _3316_ _0484_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6827_ _2824_ _2820_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6758_ _2799_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__inv_2
X_6689_ _2765_ _2885_ _2803_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__o21ai_1
X_5709_ _0353_ egd_top.BitStream_buffer.BS_buffer\[1\] _0355_ _0947_ vssd1 vssd1 vccd1
+ vccd1 _2042_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _3260_ _0345_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__nand2_2
X_5991_ _2315_ _2319_ _2320_ _2321_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__and4b_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942_ _1146_ _3502_ _3288_ _3505_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_59_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6612_ _2793_ _2809_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__nor2_1
X_4873_ _1211_ _1212_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3824_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _3362_ sky130_fd_sc_hd__buf_2
X_6543_ egd_top.exp_golomb_decoding.te_range\[2\] vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__inv_2
X_3755_ _3292_ _3219_ vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__and2_1
X_3686_ egd_top.BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__clkbuf_4
X_6474_ _2701_ _2700_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5425_ _0822_ _3368_ _1759_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5356_ _0420_ _0439_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4307_ _3295_ _3246_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__nand2_1
X_5287_ _3295_ _3306_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__nand2_1
X_4238_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__clkbuf_2
X_7026_ _3072_ _3073_ clknet_1_1__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4169_ _0512_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3540_ net35 _3098_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5210_ _1502_ _1517_ _1531_ _1546_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__and4_1
X_6190_ _2492_ _2504_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__and2_1
X_5141_ _1350_ _0621_ _1478_ _0624_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__o22ai_1
X_5072_ _0697_ _3490_ _3483_ _3493_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ _0366_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5974_ _0455_ _0733_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4925_ _3427_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _1264_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4856_ egd_top.BitStream_buffer.BS_buffer\[84\] _0494_ _0496_ _1192_ _1195_ vssd1
+ vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__a221oi_1
X_3807_ _3234_ _3323_ vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6526_ _2731_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4787_ _3427_ _3358_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__nand2_1
X_3738_ egd_top.BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6457_ net1 _0733_ net43 vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__mux2_1
X_3669_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__buf_2
X_5408_ _3263_ _3395_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6388_ _2640_ _2624_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and2_1
X_5339_ _0354_ egd_top.BitStream_buffer.BS_buffer\[126\] _0356_ egd_top.BitStream_buffer.BS_buffer\[127\]
+ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__a22o_1
X_7009_ _3066_ _3067_ clknet_1_1__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_0__3068_ _3068_ vssd1 vssd1 vccd1 vccd1 clknet_0__3068_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4710_ _1036_ _1042_ _1046_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__and4_1
X_5690_ _3344_ _3451_ _3354_ _3455_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__a221oi_1
X_4641_ _0980_ _0981_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4572_ egd_top.BitStream_buffer.BS_buffer\[82\] _0494_ _0496_ egd_top.BitStream_buffer.BS_buffer\[83\]
+ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__a221oi_1
X_3523_ _3082_ _3083_ _3084_ vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__o21ai_1
X_6311_ net6 _3372_ _2470_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__mux2_1
X_6242_ _2540_ _2536_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__and2_1
X_6173_ _2493_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
X_5124_ egd_top.BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__inv_2
X_5055_ _3414_ _3401_ _3418_ _3405_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4006_ _3234_ _0345_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5957_ _0383_ _0366_ _2287_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__o21ai_1
X_4908_ _0607_ _3326_ _0593_ _3330_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5888_ _2210_ _2214_ _2217_ _2219_ vssd1 vssd1 vccd1 vccd1 _2220_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4839_ _1175_ _0427_ _1176_ _1177_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6509_ net16 _0510_ _2707_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__3031_ clknet_0__3031_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3031_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6860_ _3033_ _3034_ clknet_1_1__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6791_ _2954_ _2900_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__nand2_1
X_5811_ _3462_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _2143_
+ sky130_fd_sc_hd__nand2_1
X_5742_ _2073_ _2074_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5673_ _3327_ _3360_ _3336_ _3364_ _2005_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__a221oi_1
X_4624_ _0814_ _3314_ _0964_ _3318_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4555_ _0892_ _0427_ _0893_ _0895_ _0896_ vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4486_ _3371_ _3362_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__nand2_1
X_6225_ net16 _3213_ _2516_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__mux2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _2481_ _3197_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__and2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5107_ _0471_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1445_
+ sky130_fd_sc_hd__nand2_1
X_6087_ _0411_ _3192_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__nand2_1
X_5038_ _1346_ _3332_ _1375_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__o21ai_1
X_6989_ _3063_ _3064_ clknet_1_1__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 la_data_out_18_16[0] sky130_fd_sc_hd__buf_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4340_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__buf_2
X_4271_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__clkbuf_4
X_6010_ _2331_ _2335_ _2338_ _2340_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6912_ _3045_ _3046_ clknet_1_0__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6843_ clknet_1_0__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6774_ _2966_ _2864_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3986_ _0328_ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5725_ _0433_ _3163_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__nand2_1
X_5656_ _3269_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _1989_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4607_ _0872_ _0946_ _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__nand3_1
XFILLER_0_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5587_ _3205_ _0347_ _1919_ _1920_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__a211oi_1
X_4538_ _3174_ _0361_ _3177_ _0364_ _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__a221oi_1
X_4469_ _3295_ _3238_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__nand2_1
X_6208_ _2517_ _2513_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__and2_1
X_7188_ _0138_ _0299_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[126\]
+ sky130_fd_sc_hd__dfxtp_1
X_6139_ net47 _3124_ _3125_ _3156_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__or4b_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3840_ _3377_ vssd1 vssd1 vccd1 vccd1 _3378_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3771_ _3308_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5510_ _0583_ _0510_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6490_ _2706_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ _3459_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _1776_
+ sky130_fd_sc_hd__nand2_1
X_5372_ _1706_ _1707_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7111_ _0061_ _0222_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_4323_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__inv_2
X_7042_ _3075_ _3076_ clknet_1_1__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__o21ai_2
X_4254_ _3292_ _0553_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__and2_1
X_4185_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6826_ _3015_ _3016_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6757_ _2948_ _2950_ vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3969_ _3251_ _3470_ vssd1 vssd1 vccd1 vccd1 _3507_ sky130_fd_sc_hd__and2_2
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5708_ _1026_ _0350_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6688_ _2764_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1
+ vccd1 vccd1 _2885_ sky130_fd_sc_hd__and2_1
X_5639_ _0589_ _0595_ _0584_ _0599_ _1972_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__3065_ clknet_0__3065_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3065_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5990_ _0513_ _0746_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__nand2_1
X_4941_ _3483_ _3490_ _0693_ _3493_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4872_ _0588_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _1212_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6611_ _2773_ _2774_ _2783_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__nand3_4
X_3823_ _3360_ vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__buf_2
XFILLER_0_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3754_ _3277_ _3116_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__nor2_4
X_6542_ net25 _2742_ net24 vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__and3b_1
XFILLER_0_27_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3685_ _3222_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__buf_2
X_6473_ _2699_ egd_top.BitStream_buffer.pc_previous\[4\] egd_top.BitStream_buffer.pc_previous\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5424_ _3371_ _3376_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5355_ _0434_ _0418_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__nand2_1
X_5286_ _3395_ _3254_ _3402_ _3258_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__a221oi_1
X_4306_ egd_top.BitStream_buffer.BS_buffer\[19\] vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4237_ _3260_ _0552_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__and2_1
X_7025_ clknet_1_0__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__buf_1
XFILLER_0_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4168_ _3226_ _0483_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__and2_1
X_4099_ _3278_ _0407_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6809_ _2989_ _3000_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5140_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__inv_2
X_5071_ _3496_ _0329_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nand2_1
X_4022_ _3278_ _0345_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5973_ _0450_ _3152_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4924_ _3453_ _3401_ _3414_ _3405_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4855_ _1193_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4786_ _3449_ _3401_ _3453_ _3405_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__a221oi_1
X_3806_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__clkbuf_4
X_3737_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__clkbuf_4
X_6525_ _2730_ _3080_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6456_ _2687_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
X_3668_ _3207_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
X_5407_ _3255_ _3223_ _3432_ _3229_ _1741_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__a221oi_2
X_3599_ net34 net33 vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__or2_1
X_6387_ net13 _0927_ _2620_ vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__mux2_1
X_5338_ _0383_ _0351_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__nor2_1
X_7008_ _3066_ _3067_ clknet_1_1__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__o21ai_2
X_5269_ _1478_ _0621_ _1605_ _0624_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _3390_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _0981_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4571_ _0911_ _0912_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6310_ _2587_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
X_3522_ net38 vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__inv_2
X_6241_ net11 _3306_ _2515_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__mux2_1
X_6172_ _2491_ _2492_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__and2_1
X_5123_ _0442_ _0521_ _0448_ _0525_ _1460_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__a221oi_1
X_5054_ _1261_ _3408_ _1391_ _3411_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__o22ai_1
X_4005_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5956_ _0369_ _3205_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__nand2_1
X_5887_ _0510_ _0613_ _0515_ _0617_ _2218_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__a221oi_1
X_4907_ _1215_ _3332_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4838_ _0892_ _0439_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4769_ _1078_ _3332_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6508_ _2719_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
X_6439_ net13 _1039_ _2656_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold10 egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__3030_ clknet_0__3030_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3030_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6790_ _2980_ _2869_ _2982_ vssd1 vssd1 vccd1 vccd1 _2983_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5810_ _3458_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _2142_
+ sky130_fd_sc_hd__nand2_1
X_5741_ _0502_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _2074_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5672_ _1111_ _3367_ _2004_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4623_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4554_ _0425_ _0439_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6224_ _2528_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4485_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__inv_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ net7 _0634_ _2480_ vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__mux2_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5106_ _0435_ _0445_ _0447_ _0741_ _1443_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__a221oi_1
X_6086_ _2407_ _2410_ _2412_ _2415_ vssd1 vssd1 vccd1 vccd1 _2416_ sky130_fd_sc_hd__and4_1
X_5037_ _3335_ _0569_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6988_ _3063_ _3064_ clknet_1_0__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5939_ _0810_ _3484_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 la_data_out_18_16[1] sky130_fd_sc_hd__buf_12
XFILLER_0_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4270_ _0613_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__buf_2
X_6911_ _3045_ _3046_ clknet_1_0__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6842_ clknet_1_1__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6773_ _2954_ _2956_ vssd1 vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3985_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__clkbuf_4
X_5724_ _0429_ _0733_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5655_ _3262_ _0675_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4606_ _0633_ _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5586_ _0353_ egd_top.BitStream_buffer.BS_buffer\[0\] _0355_ _0796_ vssd1 vssd1 vccd1
+ vccd1 _1920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4537_ _0877_ _0367_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__o21ai_1
X_4468_ egd_top.BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__inv_2
X_6207_ net7 _3275_ _2516_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__mux2_1
X_7187_ _0137_ _0298_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[127\]
+ sky130_fd_sc_hd__dfxtp_1
X_6138_ _2347_ _2467_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__nor2_1
X_4399_ _0434_ _0741_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__nand2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _0327_ egd_top.BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _2399_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3770_ _3307_ _3220_ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5440_ _0836_ _3435_ _3438_ _3449_ _1774_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5371_ _0503_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _1707_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7110_ _0060_ _0221_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_4322_ _3344_ _3343_ _3354_ _3347_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7041_ _3075_ _3076_ clknet_1_1__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__o21ai_2
X_4253_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__clkbuf_4
X_4184_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__buf_2
XFILLER_0_89_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6825_ _3011_ vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__inv_2
X_3968_ _3500_ _3502_ _3503_ _3505_ vssd1 vssd1 vccd1 vccd1 _3506_ sky130_fd_sc_hd__o22ai_1
X_6756_ _2760_ _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__nor2_1
X_5707_ _1997_ _2011_ _2024_ _2039_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6687_ _2882_ _2883_ _2801_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3899_ _3436_ vssd1 vssd1 vccd1 vccd1 _3437_ sky130_fd_sc_hd__clkbuf_2
X_5638_ _0790_ _0602_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__o21ai_1
X_5569_ _3474_ _3275_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4940_ _3496_ _0339_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4871_ _0583_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _1211_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6610_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1 vccd1 vccd1
+ _2808_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3822_ _3359_ vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__clkbuf_2
X_6541_ _2741_ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__inv_2
X_3753_ _3290_ vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3684_ _3221_ vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__clkbuf_2
X_6472_ _3120_ _3090_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5423_ _3327_ _3343_ _3336_ _3347_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5354_ _0430_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1690_
+ sky130_fd_sc_hd__nand2_1
X_4305_ egd_top.BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__clkbuf_4
X_5285_ _1619_ _1620_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4236_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__clkbuf_4
X_7024_ _3026_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__buf_4
X_4167_ _0509_ _0510_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4098_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6808_ _2999_ vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__inv_2
X_6739_ _2930_ _2933_ _2934_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__3047_ clknet_0__3047_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3047_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _1141_ _3472_ _1405_ _1406_ _1407_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__o2111a_1
X_4021_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _1161_ _0426_ _2300_ _2301_ _2302_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__o2111a_1
X_4923_ _1124_ _3408_ _1261_ _3411_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__o22ai_1
X_4854_ _0503_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _1194_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4785_ _0985_ _3408_ _1124_ _3411_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3805_ _3342_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__buf_2
X_3736_ _3250_ _3254_ _3255_ _3258_ _3273_ vssd1 vssd1 vccd1 vccd1 _3274_ sky130_fd_sc_hd__a221oi_2
X_6524_ net11 _0522_ _2706_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6455_ _2686_ _2668_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3667_ _3206_ _3197_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__and2_1
X_5406_ _1739_ _1740_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__nand2_1
X_6386_ _2639_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
X_3598_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__buf_2
X_5337_ _1629_ _1643_ _1657_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__and4_1
X_5268_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__inv_2
X_7007_ _3066_ _3067_ clknet_1_0__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__o21ai_2
X_4219_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__buf_2
X_5199_ _3496_ _0334_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4570_ _0503_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0912_
+ sky130_fd_sc_hd__nand2_1
X_3521_ net36 net35 vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6240_ _2539_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
X_6171_ _3165_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__buf_8
X_5122_ _0772_ _0528_ _0923_ _0531_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__o22ai_1
X_5053_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__inv_2
X_4004_ _0347_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5955_ _0796_ _0347_ _2284_ _2285_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5886_ _2096_ _0620_ _0481_ _0623_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__o22ai_1
X_4906_ _3335_ _0597_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__nand2_1
X_4837_ _0434_ _0461_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4768_ _3335_ _0593_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__nand2_1
X_3719_ _3256_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__clkbuf_2
X_6507_ _2718_ _2689_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__and2_1
X_4699_ _0434_ _1039_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__nand2_1
X_6438_ _2675_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
X_6369_ net4 _0597_ _2620_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5740_ _0498_ _0534_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5671_ _3370_ _3322_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__nand2_1
X_4622_ _3296_ _3281_ _3286_ _3246_ _0962_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__a221oi_1
X_4553_ _0434_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4484_ _3354_ _3343_ _0662_ _3347_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__a221oi_1
X_6223_ _2513_ _2527_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__and2_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _2479_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__clkbuf_4
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _1441_ _1442_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__nand2_1
X_6085_ _3476_ _0389_ _3482_ _0392_ _2414_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__a221oi_1
X_5036_ _1363_ _1367_ _1370_ _1373_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__and4_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6987_ _3063_ _3064_ clknet_1_0__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__o21ai_2
X_5938_ _3479_ _3287_ vssd1 vssd1 vccd1 vccd1 _2269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5869_ _2194_ _2198_ _2199_ _2200_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__and4b_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 la_data_out_18_16[2] sky130_fd_sc_hd__buf_12
XFILLER_0_39_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6910_ _3045_ _3046_ clknet_1_0__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__o21ai_2
X_6841_ _3029_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__buf_1
X_3984_ _0327_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__clkbuf_4
X_6772_ _2958_ _2955_ _2865_ vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5723_ _1291_ _0408_ _2053_ _2054_ _2055_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__o2111a_1
X_5654_ _3439_ _3222_ _0683_ _3228_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4605_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__clkbuf_4
X_5585_ _0881_ _0350_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4536_ _0370_ _3171_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__nand2_1
X_4467_ _3432_ _3254_ _3439_ _3258_ _0808_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a221oi_1
X_6206_ _2515_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__clkbuf_4
X_7186_ _0136_ _0297_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_4398_ egd_top.BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__clkbuf_4
X_6137_ _3149_ _2466_ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__nor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _0322_ _0801_ vssd1 vssd1 vccd1 vccd1 _2398_ sky130_fd_sc_hd__nand2_1
X_5019_ _3212_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _0499_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _1706_
+ sky130_fd_sc_hd__nand2_1
X_4321_ _0661_ _3350_ _0663_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__o21ai_1
X_7040_ _3075_ _3076_ clknet_1_1__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__o21ai_2
X_4252_ _0595_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4183_ _3312_ _0484_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nand2_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6824_ _3014_ _2966_ vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__nand2_1
X_3967_ _3504_ vssd1 vssd1 vccd1 vccd1 _3505_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6755_ _2914_ vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5706_ _2028_ _2030_ _2033_ _2038_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__and4_1
X_6686_ _2848_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] vssd1 vssd1 vccd1
+ vccd1 _2883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3898_ _3283_ _3398_ vssd1 vssd1 vccd1 vccd1 _3436_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5637_ _0605_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _1971_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5568_ _1891_ _1894_ _1897_ _1901_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__and4_1
X_4519_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__inv_2
X_5499_ _0514_ _0442_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__nand2_1
X_7169_ _0119_ _0280_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4870_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3821_ _3289_ _3323_ vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__and2_1
X_6540_ net18 net17 vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__nand2_1
X_3752_ _3289_ _3220_ vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3683_ _3217_ _3220_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__and2_1
X_6471_ egd_top.BitStream_buffer.pc_previous\[6\] _2700_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[6\]
+ sky130_fd_sc_hd__xor2_4
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5422_ _0601_ _3350_ _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5353_ _0873_ _0409_ _1686_ _1687_ _1688_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__o2111a_1
X_4304_ _3255_ _3254_ _3432_ _3258_ _0646_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _3270_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _1620_
+ sky130_fd_sc_hd__nand2_1
X_4235_ _0578_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__clkbuf_2
X_7023_ _3023_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__buf_4
X_4166_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4097_ _0425_ _0427_ _0431_ _0436_ _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_77_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6807_ _2998_ _2825_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4999_ _0563_ _0611_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6738_ net24 net25 vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6669_ _2866_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4020_ _0363_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5971_ _0877_ _0438_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__or2_1
X_4922_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4853_ _0499_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _1193_
+ sky130_fd_sc_hd__nand2_1
X_4784_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3804_ _3341_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__clkbuf_2
X_3735_ _3265_ _3272_ vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__nand2_1
X_6523_ _2729_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6454_ net8 _0418_ net43 vssd1 vssd1 vccd1 vccd1 _2686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ _3245_ _3264_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3666_ net8 _3205_ _3158_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3597_ _3151_ _3141_ _3081_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__o21ai_1
X_6385_ _2638_ _2624_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__and2_1
X_5336_ _1661_ _1663_ _1666_ _1671_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__and4_1
X_5267_ _0927_ _0596_ _0611_ _0600_ _1603_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__a221oi_1
X_7006_ _3066_ _3067_ clknet_1_0__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__o21ai_2
X_4218_ _0561_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__clkbuf_2
X_5198_ _3500_ _3472_ _1532_ _1533_ _1534_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__o2111a_1
Xclkbuf_0__3065_ _3065_ vssd1 vssd1 vccd1 vccd1 clknet_0__3065_ sky130_fd_sc_hd__clkbuf_16
X_4149_ _0492_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3520_ net37 vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__inv_2
X_6170_ net2 _0695_ _2480_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__mux2_1
X_5121_ _1452_ _1456_ _1457_ _1458_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__and4b_1
XFILLER_0_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _1377_ _1381_ _1385_ _1389_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4003_ _0346_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5954_ _0353_ _3497_ _0355_ _0701_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4905_ _1232_ _1236_ _1240_ _1243_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__and4_1
X_5885_ _0573_ _0595_ _0577_ _0599_ _2216_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__a221oi_1
X_4836_ _0430_ _0894_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__nand2_1
X_4767_ _1095_ _1099_ _1103_ _1106_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__and4_1
X_6506_ net2 _1192_ _2707_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3718_ _3119_ _3220_ vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__and2_1
X_4698_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6437_ _2674_ _2668_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__and2_1
X_3649_ net12 _3192_ _3158_ vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__mux2_1
X_6368_ _2627_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5319_ _1653_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__nand2_1
X_6299_ net39 vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5670_ _0657_ _3342_ _0818_ _3346_ _2002_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _0960_ _3291_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4552_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__clkbuf_4
X_4483_ _0822_ _3350_ _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__o21ai_1
X_6222_ net2 _3238_ _2516_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6153_ _2471_ _3133_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__nand2_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _0855_ _0395_ _2413_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__o21ai_1
X_5104_ _0456_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _1442_
+ sky130_fd_sc_hd__nand2_1
X_5035_ _3432_ _3305_ _3439_ _3310_ _1372_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__a221oi_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6986_ clknet_1_1__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__buf_1
X_5937_ _3474_ _3296_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5868_ _0513_ _0452_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5799_ _2129_ _2130_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__nand2_1
X_4819_ _0354_ egd_top.BitStream_buffer.BS_buffer\[122\] _0356_ _3195_ vssd1 vssd1
+ vccd1 vccd1 _1159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[0] sky130_fd_sc_hd__buf_12
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[0] sky130_fd_sc_hd__buf_12
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6840_ wb_clk_i _3026_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__or2b_2
X_6771_ _2963_ _2964_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__nand2_1
X_3983_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5722_ _1018_ _0421_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5653_ _1984_ _1985_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4604_ _0907_ _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__nor2_1
X_5584_ _1875_ _1889_ _1902_ _1917_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4535_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4466_ _0806_ _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7185_ _0135_ _0296_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_6205_ _2471_ _3132_ _2474_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__nand3_4
X_4397_ _0430_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__nand2_1
X_6136_ _2404_ _2464_ _2465_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__nand3_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _2395_ _2396_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__nor2_1
X_5018_ _1290_ _1355_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__nand3_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6969_ _3057_ _3058_ clknet_1_0__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4320_ _3353_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__nand2_1
X_4251_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4182_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6823_ _2998_ _2978_ _2861_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3966_ _3260_ _3470_ vssd1 vssd1 vccd1 vccd1 _3504_ sky130_fd_sc_hd__nand2_2
X_6754_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _2914_ vssd1 vssd1 vccd1
+ vccd1 _2948_ sky130_fd_sc_hd__nor2_1
X_5705_ _2034_ _2035_ _2036_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6685_ _2847_ _2760_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3897_ _3434_ vssd1 vssd1 vccd1 vccd1 _3435_ sky130_fd_sc_hd__buf_2
X_5636_ _0765_ _0575_ _0916_ _0579_ _1969_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_5_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5567_ _3340_ _3451_ _3344_ _3455_ _1900_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5498_ _0509_ _0538_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__nand2_1
X_4518_ _0858_ _3490_ _0700_ _3493_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__o221a_1
X_4449_ _0615_ _0614_ _0589_ _0618_ _0791_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__a221oi_1
X_7168_ _0118_ _0279_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6119_ _0562_ _1210_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__nand2_1
X_7099_ _0049_ _0210_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3062_ clknet_0__3062_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3062_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3820_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__buf_2
X_3751_ _3277_ _3214_ vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__nor2_4
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3682_ _3219_ vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__buf_2
X_6470_ _2699_ egd_top.BitStream_buffer.pc_previous\[4\] egd_top.BitStream_buffer.pc_previous\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__and3_2
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5421_ _3353_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _1756_
+ sky130_fd_sc_hd__nand2_1
X_5352_ _0349_ _0422_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__or2_1
X_4303_ _0644_ _0645_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nand2_1
X_5283_ _3263_ _1130_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__nand2_1
X_7022_ _3069_ _3070_ clknet_1_1__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__o21ai_2
X_4234_ _3119_ _0553_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4165_ _0508_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4096_ _0437_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6806_ _2990_ _2997_ vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__nor2_1
X_4998_ _1331_ _1333_ _1336_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6737_ _2932_ _2900_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3949_ _3468_ _3472_ _3477_ _3481_ _3486_ vssd1 vssd1 vccd1 vccd1 _3487_ sky130_fd_sc_hd__o2111a_1
X_6668_ _2860_ _2861_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__nand2_1
X_6599_ _2796_ _2767_ _2780_ _2791_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__o211ai_4
X_5619_ _1951_ _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _0433_ _3171_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__nand2_1
X_4921_ _1247_ _1251_ _1255_ _1259_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__and4_1
X_4852_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__clkbuf_4
X_3803_ _3242_ _3323_ vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4783_ _1110_ _1114_ _1118_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__and4_1
X_3734_ _3270_ _3271_ vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__nand2_1
X_6522_ _2728_ _3080_ vssd1 vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__and2_1
X_6453_ _2685_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
X_3665_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__buf_2
X_5404_ _3237_ _3250_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3596_ _3150_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__clkbuf_4
X_6384_ net14 _0776_ _2620_ vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__mux2_1
X_5335_ _1667_ _1668_ _1669_ _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__and4_1
X_5266_ _1601_ _0603_ _1602_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7005_ _3066_ _3067_ clknet_1_0__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__o21ai_2
X_4217_ _3234_ _0552_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__and2_1
X_5197_ _0704_ _3485_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__or2_1
X_4148_ _3278_ _0483_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _0420_ _0422_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5120_ _0514_ _0919_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__nand2_1
X_5051_ _0818_ _3379_ _0607_ _3383_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__a221oi_1
X_4002_ _3242_ _0345_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _3488_ _0350_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__nor2_1
X_4904_ _3255_ _3305_ _3432_ _3310_ _1242_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5884_ _1082_ _0602_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__o21ai_1
X_4835_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__inv_2
X_4766_ _3250_ _3305_ _3255_ _3310_ _1105_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3717_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__clkbuf_4
X_6505_ _2717_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4697_ _0430_ _0741_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__nand2_1
X_6436_ net14 _0894_ _2656_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__mux2_1
X_3648_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6367_ _2626_ _2624_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__and2_1
X_3579_ egd_top.BitStream_buffer.pc_previous\[6\] _3120_ vssd1 vssd1 vccd1 vccd1 _3137_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5318_ _3463_ egd_top.BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _1654_
+ sky130_fd_sc_hd__nand2_1
X_6298_ net9 _3418_ _2550_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__mux2_1
X_5249_ _1579_ _1583_ _1584_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__and4b_1
Xclkbuf_0__3047_ _3047_ vssd1 vssd1 vccd1 vccd1 clknet_0__3047_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4620_ _3295_ _3213_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4551_ _0430_ _0435_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__nand2_1
X_4482_ _3353_ _0823_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nand2_1
X_6221_ _2526_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _2477_ _2478_ _3089_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a21oi_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _0451_ _1039_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__nand2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _0398_ _0339_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__nand2_1
X_5034_ _1241_ _3314_ _1371_ _3318_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__o22ai_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6985_ _3026_ vssd1 vssd1 vccd1 vccd1 _3064_ sky130_fd_sc_hd__buf_4
X_5936_ _2256_ _2259_ _2262_ _2266_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__and4_1
XFILLER_0_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5867_ _0508_ _0457_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5798_ _3389_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _2130_
+ sky130_fd_sc_hd__nand2_1
X_4818_ _1157_ _0351_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4749_ _3212_ _1089_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[1] sky130_fd_sc_hd__buf_12
X_6419_ _2662_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[1] sky130_fd_sc_hd__buf_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3982_ _3316_ _3469_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__and2_1
X_6770_ _2924_ _2900_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__nand2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5721_ _0416_ _3189_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nand2_1
X_5652_ _3244_ _3255_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5583_ _1906_ _1908_ _1911_ _1916_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__and4_1
X_4603_ _0926_ _0944_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4534_ _3180_ _0348_ _0874_ _0875_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4465_ _3270_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _0807_
+ sky130_fd_sc_hd__nand2_1
X_7184_ _0134_ _0295_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4396_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__clkbuf_4
X_6204_ _2514_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _0632_ _3509_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__nand2_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _3507_ egd_top.BitStream_buffer.BS_buffer\[28\] _3510_ egd_top.BitStream_buffer.BS_buffer\[29\]
+ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__a22o_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5017_ _0633_ _0695_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6968_ _3057_ _3058_ clknet_1_0__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6899_ _3042_ _3043_ clknet_1_1__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__o21ai_2
X_5919_ _3385_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _2250_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _3289_ _0553_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__and2_1
X_4181_ _0524_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6822_ _3012_ _2865_ vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6753_ _2763_ _2920_ vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _3503_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5704_ _0337_ egd_top.BitStream_buffer.BS_buffer\[19\] vssd1 vssd1 vccd1 vccd1 _2037_
+ sky130_fd_sc_hd__nand2_1
X_6684_ _2876_ _2880_ _2818_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__nand3_1
X_3896_ _3433_ vssd1 vssd1 vccd1 vccd1 _3434_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5635_ _1967_ _1968_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5566_ _1898_ _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__nand2_1
X_5497_ _0916_ _0494_ _0496_ _0518_ _1831_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__a221oi_1
X_4517_ _3496_ _0695_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__nand2_1
X_4448_ _0622_ _0621_ _0790_ _0624_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__o22ai_1
X_4379_ _0720_ _0367_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__o21ai_1
X_7167_ _0117_ _0278_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_6118_ _2443_ _2445_ _2447_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__and3_1
X_7098_ _0048_ _0209_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _1378_ _3423_ _2378_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3750_ egd_top.BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3681_ _3120_ _3218_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _3219_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5420_ _0564_ _3326_ _0551_ _3330_ _1754_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5351_ _0417_ _3180_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__nand2_1
X_5282_ _3250_ _3223_ _3255_ _3229_ _1617_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__a221oi_1
X_4302_ _3270_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _0645_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4233_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__clkbuf_4
X_7021_ _3069_ _3070_ clknet_1_1__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__o21ai_2
X_4164_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4095_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6805_ _2995_ _2996_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__nand2_1
X_6736_ _2931_ vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__inv_2
X_4997_ _0452_ _0537_ _0746_ _0541_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__a221oi_1
X_3948_ _3483_ _3485_ vssd1 vssd1 vccd1 vccd1 _3486_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6667_ _2864_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__inv_4
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3879_ _3416_ vssd1 vssd1 vccd1 vccd1 _3417_ sky130_fd_sc_hd__buf_2
X_6598_ _2760_ _2758_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__nand2_1
X_5618_ _0502_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _1952_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5549_ _0971_ _3367_ _1882_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__3044_ clknet_0__3044_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3044_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4920_ _0657_ _3379_ _0818_ _3383_ _1258_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__a221oi_1
X_4851_ _0529_ _0486_ _1190_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3802_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__buf_2
XFILLER_0_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4782_ _3336_ _3379_ _0657_ _3383_ _1121_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3733_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__clkbuf_4
X_6521_ net12 _0518_ _2706_ vssd1 vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6452_ _2684_ _2668_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__and2_1
X_3664_ _3204_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_1
X_5403_ _3150_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__o21ai_1
X_3595_ _3149_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__inv_2
X_6383_ _2637_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
X_5334_ _0338_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1670_
+ sky130_fd_sc_hd__nand2_1
X_5265_ _0606_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _1602_
+ sky130_fd_sc_hd__nand2_1
X_5196_ _3480_ _0324_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__nand2_1
X_7004_ _3066_ _3067_ clknet_1_1__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__o21ai_2
X_4216_ _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4147_ _0481_ _0486_ _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__o21ai_1
X_4078_ _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6719_ _2758_ _2788_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5050_ _1386_ _1387_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__nand2_1
X_4001_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5952_ _2240_ _2254_ _2267_ _2282_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4903_ _1104_ _3314_ _1241_ _3318_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5883_ _0605_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _2215_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4834_ _1022_ _0409_ _1171_ _1172_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4765_ _0964_ _3314_ _1104_ _3318_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o22ai_1
X_3716_ _3253_ vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__buf_2
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6504_ _2716_ _2689_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__and2_1
X_4696_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__inv_2
X_6435_ _2673_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
X_3647_ _3191_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
X_3578_ egd_top.BitStream_buffer.pc\[6\] _3123_ _3135_ vssd1 vssd1 vccd1 vccd1 _3136_
+ sky130_fd_sc_hd__or3b_1
X_6366_ net5 _0593_ _2620_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__mux2_1
X_5317_ _3459_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _1653_
+ sky130_fd_sc_hd__nand2_1
X_6297_ _2578_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
X_5248_ _0514_ _0534_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__nand2_1
X_5179_ _0607_ _3379_ _0593_ _3383_ _1515_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4481_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__clkbuf_4
X_6220_ _2525_ _2513_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__and2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _2471_ _3125_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__nand2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _0420_ _0427_ _1437_ _1438_ _1439_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__o2111a_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _0708_ _0375_ _0865_ _0378_ _2411_ vssd1 vssd1 vccd1 vccd1 _2412_ sky130_fd_sc_hd__a221oi_1
X_5033_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__inv_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6984_ _3023_ vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5935_ _0662_ _3451_ _0823_ _3455_ _2265_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5866_ _0768_ _0493_ _0495_ _0919_ _2197_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__a221oi_1
X_4817_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5797_ _3385_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _2129_
+ sky130_fd_sc_hd__nand2_1
X_4748_ _1017_ _1087_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__nand3_2
X_4679_ _0354_ egd_top.BitStream_buffer.BS_buffer\[121\] _0356_ egd_top.BitStream_buffer.BS_buffer\[122\]
+ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__a22o_1
X_6418_ _2661_ _2645_ vssd1 vssd1 vccd1 vccd1 _2662_ sky130_fd_sc_hd__and2_1
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[2] sky130_fd_sc_hd__buf_12
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[2] sky130_fd_sc_hd__buf_12
X_6349_ _2613_ _2601_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__and2_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3981_ _0323_ _0324_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__nand2_1
X_5720_ _0411_ _3183_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _3236_ _3432_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5582_ _1912_ _1913_ _1914_ _1915_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602_ _0931_ _0936_ _0940_ _0943_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__and4_1
X_4533_ _0354_ egd_top.BitStream_buffer.BS_buffer\[120\] _0356_ egd_top.BitStream_buffer.BS_buffer\[121\]
+ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _3263_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _0806_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6203_ _2512_ _2513_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7183_ _0133_ _0294_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ sky130_fd_sc_hd__dfxtp_2
X_4395_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__inv_2
X_6134_ _2434_ _2463_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__nor2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _0653_ _3501_ _0814_ _3504_ vssd1 vssd1 vccd1 vccd1 _2395_ sky130_fd_sc_hd__o22ai_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5016_ _1322_ _1354_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__nor2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _3057_ _3058_ clknet_1_1__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__o21ai_2
X_5918_ _0657_ _3360_ _0818_ _3364_ _2248_ vssd1 vssd1 vccd1 vccd1 _2249_ sky130_fd_sc_hd__a221oi_1
X_6898_ _3042_ _3043_ clknet_1_1__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5849_ _0720_ _0438_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4180_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6821_ _3008_ _3011_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ _3501_ vssd1 vssd1 vccd1 vccd1 _3502_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6752_ _2920_ _2763_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5703_ _0332_ egd_top.BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _2036_
+ sky130_fd_sc_hd__nand2_1
X_6683_ _2817_ _2879_ _2831_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__nand3_1
X_3895_ _3278_ _3397_ vssd1 vssd1 vccd1 vccd1 _3433_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5634_ _0587_ _0510_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5565_ _3462_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _1899_
+ sky130_fd_sc_hd__nand2_1
X_5496_ _1829_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__nand2_1
X_4516_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__inv_2
X_4447_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__inv_2
X_7166_ _0116_ _0277_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_6117_ _0413_ _0536_ _0731_ _0540_ _2446_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__a221oi_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ _0370_ _3168_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__nand2_1
X_7097_ _0047_ _0208_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _3426_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _2378_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__inv_2
X_5350_ _0412_ _3174_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__nand2_1
X_5281_ _1615_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__nand2_1
X_4301_ _3263_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _0644_
+ sky130_fd_sc_hd__nand2_1
X_4232_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__clkbuf_4
X_7020_ _3069_ _3070_ clknet_1_1__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__o21ai_2
X_4163_ _3217_ _0484_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__and2_1
X_4094_ _3234_ _0407_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__nand2_1
X_6804_ _2943_ _2991_ _2993_ vssd1 vssd1 vccd1 vccd1 _2996_ sky130_fd_sc_hd__nand3_1
X_4996_ _1202_ _0544_ _1334_ _0547_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__o22ai_1
X_3947_ _3484_ vssd1 vssd1 vccd1 vccd1 _3485_ sky130_fd_sc_hd__clkbuf_2
X_6735_ _2895_ _2861_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6666_ _2820_ _2861_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__nand2_2
X_3878_ _3415_ vssd1 vssd1 vccd1 vccd1 _3416_ sky130_fd_sc_hd__clkbuf_2
X_5617_ _0498_ _0919_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__nand2_1
X_6597_ _2795_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ sky130_fd_sc_hd__inv_2
X_5548_ _3370_ _3380_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__nand2_1
X_5479_ _0434_ _0733_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__nand2_1
X_7149_ _0099_ _0260_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _0489_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _1190_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3801_ _3322_ _3326_ _3327_ _3330_ _3338_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__a221oi_1
X_6520_ _2727_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _1119_ _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3732_ _3269_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6451_ net9 _0731_ net43 vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__mux2_1
X_3663_ _3203_ _3197_ vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5402_ _1614_ _1737_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__nor2_1
X_6382_ _2636_ _2624_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5333_ _0333_ _0648_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__nand2_1
X_3594_ egd_top.BitStream_buffer.BitStream_buffer_valid_n vssd1 vssd1 vccd1 vccd1
+ _3149_ sky130_fd_sc_hd__buf_6
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5264_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5195_ _3475_ _0865_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__nand2_1
X_7003_ _3066_ _3067_ clknet_1_0__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__o21ai_2
X_4215_ _0558_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3062_ _3062_ vssd1 vssd1 vccd1 vccd1 clknet_0__3062_ sky130_fd_sc_hd__clkbuf_16
X_4146_ _0489_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0490_
+ sky130_fd_sc_hd__nand2_1
X_4077_ _3260_ _0407_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4979_ _0475_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _1318_
+ sky130_fd_sc_hd__nand2_1
X_6718_ _2787_ _2848_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6649_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4000_ egd_top.BitStream_buffer.pc\[6\] egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__and3_2
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5951_ _2271_ _2273_ _2276_ _2281_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__and4_1
X_4902_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ _0518_ _0575_ _0522_ _0579_ _2213_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__a221oi_1
X_4833_ _0720_ _0422_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4764_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ _3252_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__clkbuf_2
X_6503_ net3 _1055_ _2707_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6434_ _2672_ _2668_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__and2_1
X_4695_ _0877_ _0409_ _1033_ _1034_ _1035_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3646_ _3190_ _3166_ vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ _2625_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
X_3577_ _3134_ egd_top.BitStream_buffer.pc_previous\[4\] egd_top.BitStream_buffer.pc_previous\[5\]
+ egd_top.BitStream_buffer.pc_previous\[6\] vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__a31o_1
X_6296_ _2577_ _2559_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__and2_1
X_5316_ _0675_ _3435_ _3438_ _0836_ _1651_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__a221oi_1
X_5247_ _0509_ _0919_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__nand2_1
X_5178_ _1513_ _1514_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__nand2_1
X_4129_ _3312_ _0406_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4480_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__inv_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _3125_ _2471_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__or2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _1175_ _0439_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__or2_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _1002_ _0381_ _1141_ _0384_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__o22ai_1
X_5032_ _3213_ _3281_ _3286_ _3224_ _1369_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__a221oi_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6983_ _3060_ _3061_ clknet_1_0__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__o21ai_2
X_5934_ _2263_ _2264_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5865_ _2195_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4816_ _1107_ _1123_ _1138_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5796_ _3336_ _3360_ _0657_ _3364_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__a221oi_1
X_4747_ _0633_ _3497_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4678_ _1018_ _0351_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__nor2_1
X_6417_ net5 _0457_ _2656_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3629_ net2 _3177_ _3159_ vssd1 vssd1 vccd1 vccd1 _3178_ sky130_fd_sc_hd__mux2_1
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 la_data_out_22_19[3] sky130_fd_sc_hd__buf_12
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[3] sky130_fd_sc_hd__buf_12
X_6348_ net9 _3327_ _2469_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__mux2_1
X_6279_ _2566_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _3150_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__o21ai_1
X_4601_ _0589_ _0614_ _0584_ _0618_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__a221oi_1
X_5581_ _0337_ egd_top.BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1 _1915_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _0873_ _0351_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__nor2_1
X_4463_ _0639_ _3223_ _0801_ _3229_ _0804_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6202_ _3165_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__buf_8
X_7182_ _0132_ _0293_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_4394_ _0365_ _0409_ _0732_ _0734_ _0736_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__3068_ clknet_0__3068_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3068_
+ sky130_fd_sc_hd__clkbuf_16
X_6133_ _2448_ _2462_ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__nand2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6064_ _1007_ _3489_ _0861_ _3492_ _2393_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__o221a_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _1337_ _1353_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__nand2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6966_ _3057_ _3058_ clknet_1_1__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__o21ai_2
X_5917_ _1378_ _3367_ _2247_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__o21ai_1
X_6897_ _3042_ _3043_ clknet_1_1__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__o21ai_2
X_5848_ _0433_ _3168_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5779_ _3269_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _2111_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6820_ _3010_ _2825_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3963_ _3267_ _3470_ vssd1 vssd1 vccd1 vccd1 _3501_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6751_ _2942_ _2944_ _2818_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__nand3_1
X_3894_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _3432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5702_ _0327_ _3246_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__nand2_1
X_6682_ _2877_ _2878_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5633_ _0582_ _0515_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__nand2_1
X_5564_ _3458_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _1898_
+ sky130_fd_sc_hd__nand2_1
X_4515_ _3483_ _3472_ _0853_ _0854_ _0856_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5495_ _0503_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _1830_
+ sky130_fd_sc_hd__nand2_1
X_4446_ _0597_ _0596_ _0569_ _0600_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__a221oi_1
X_4377_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__inv_2
X_7165_ _0115_ _0276_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_6116_ _1037_ _0543_ _1175_ _0546_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__o22ai_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _0046_ _0207_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _3340_ _3400_ _3344_ _3404_ _2376_ vssd1 vssd1 vccd1 vccd1 _2377_ sky130_fd_sc_hd__a221oi_1
X_6949_ _3054_ _3055_ clknet_1_0__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4300_ _3224_ _3223_ _0639_ _3229_ _0642_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__a221oi_1
X_5280_ _3245_ _3271_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ _0574_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__clkbuf_2
X_4162_ egd_top.BitStream_buffer.BS_buffer\[80\] _0494_ _0496_ egd_top.BitStream_buffer.BS_buffer\[81\]
+ _0505_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__a221oi_1
X_4093_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
X_6803_ _2992_ _2994_ vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__nand2_1
X_4995_ egd_top.BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__inv_2
X_3946_ _3226_ _3470_ vssd1 vssd1 vccd1 vccd1 _3484_ sky130_fd_sc_hd__nand2_1
X_6734_ _2929_ _2869_ vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6665_ _2862_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__inv_2
X_3877_ _3267_ _3398_ vssd1 vssd1 vccd1 vccd1 _3415_ sky130_fd_sc_hd__and2_1
X_5616_ _0923_ _0485_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__o21ai_1
X_6596_ _2740_ _2745_ _2794_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5547_ _3336_ _3342_ _0657_ _3346_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__a221oi_1
X_5478_ _0430_ _0731_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__nand2_1
X_4429_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__inv_2
X_7148_ _0098_ _0259_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7079_ _0029_ _0190_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _3331_ _3332_ _3337_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__o21ai_1
X_4780_ _3390_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _1120_
+ sky130_fd_sc_hd__nand2_1
X_3731_ _3268_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6450_ _2683_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3662_ net9 _3202_ _3158_ vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5401_ _3212_ _1736_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__nor2_1
X_3593_ _3147_ _3148_ _3090_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a21oi_1
X_6381_ net15 _0557_ _2620_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5332_ _0328_ _3287_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5263_ _1192_ _0576_ _0510_ _0580_ _1599_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7002_ _3066_ _3067_ clknet_1_0__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__o21ai_2
X_4214_ _3226_ _0553_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__and2_1
X_5194_ _1520_ _1523_ _1526_ _1530_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4145_ _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4978_ _0471_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _1317_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3929_ _3413_ _3431_ _3448_ _3466_ vssd1 vssd1 vccd1 vccd1 _3467_ sky130_fd_sc_hd__and4_1
X_6717_ _2907_ _2818_ _2912_ vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__nand3_1
X_6648_ _2840_ _2845_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6579_ _2768_ _2760_ _2758_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__and3_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5950_ _2277_ _2278_ _2279_ _2280_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__and4_1
X_4901_ _3238_ _3281_ _3286_ _3213_ _1239_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5881_ _2211_ _2212_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4832_ _0417_ _3168_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4763_ _3246_ _3281_ _3286_ _3238_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3714_ _3251_ _3220_ vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6502_ _2715_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4694_ _0365_ _0422_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__or2_1
X_6433_ net15 _0741_ _2656_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3645_ net13 _3189_ _3159_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__mux2_1
X_3576_ egd_top.BitStream_buffer.pc_previous\[0\] egd_top.BitStream_buffer.pc_previous\[1\]
+ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.pc_previous\[3\]
+ vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__and4_1
X_6364_ _2623_ _2624_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__and2_1
X_6295_ net10 _3414_ _2550_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__mux2_1
X_5315_ _1261_ _3442_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5246_ egd_top.BitStream_buffer.BS_buffer\[87\] _0494_ _0496_ _0765_ _1582_ vssd1
+ vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__3044_ _3044_ vssd1 vssd1 vccd1 vccd1 clknet_0__3044_ sky130_fd_sc_hd__clkbuf_16
X_5177_ _3390_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _1514_
+ sky130_fd_sc_hd__nand2_1
X_4128_ _0471_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0472_
+ sky130_fd_sc_hd__nand2_1
X_4059_ _0358_ _0373_ _0387_ _0402_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5100_ _0434_ _0413_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__nand2_1
X_6080_ _0634_ _0360_ _0796_ _0363_ _2409_ vssd1 vssd1 vccd1 vccd1 _2410_ sky130_fd_sc_hd__a221oi_1
X_5031_ _3311_ _3291_ _1368_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__o21ai_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6982_ _3060_ _3061_ clknet_1_0__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _3462_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _2264_
+ sky130_fd_sc_hd__nand2_1
X_5864_ _0502_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _2196_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ _1143_ _1145_ _1149_ _1154_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5795_ _1248_ _3367_ _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__o21ai_1
X_4746_ _1052_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__nor2_1
X_4677_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__inv_2
X_6416_ _2660_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
X_3628_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__buf_2
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[4] sky130_fd_sc_hd__buf_12
X_6347_ _2612_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3559_ _3116_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__inv_2
X_6278_ _2565_ _2559_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__and2_1
X_5229_ _1308_ _0439_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _0790_ _0621_ _0941_ _0624_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__o22ai_1
X_5580_ _0332_ egd_top.BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _1914_
+ sky130_fd_sc_hd__nand2_1
X_4531_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__inv_2
X_4462_ _0802_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6201_ net1 _3512_ _2479_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7181_ _0131_ _0292_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_4393_ _0735_ _0422_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__or2_1
X_6132_ _2452_ _2456_ _2459_ _2461_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__and4_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _3495_ _3287_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__nand2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5014_ _1341_ _1345_ _1349_ _1352_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__and4_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6965_ _3057_ _3058_ clknet_1_0__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__o21ai_2
X_5916_ _3370_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _2247_
+ sky130_fd_sc_hd__nand2_1
X_6896_ _3042_ _3043_ clknet_1_1__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5847_ _0429_ _3152_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__nand2_1
X_5778_ _3262_ _0836_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__nand2_1
X_4729_ _0568_ _0557_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6750_ _2943_ _2940_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__nand2_1
X_5701_ _0322_ _3213_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__nand2_1
X_3962_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _3500_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6681_ _2814_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1
+ vccd1 _2878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3893_ _3414_ _3417_ _3418_ _3421_ _3430_ vssd1 vssd1 vccd1 vccd1 _3431_ sky130_fd_sc_hd__a221oi_1
X_5632_ _0781_ _0555_ _0932_ _0559_ _1965_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5563_ _3449_ _3434_ _3437_ _3453_ _1896_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__a221oi_1
X_4514_ _0855_ _3485_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5494_ _0499_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _1829_
+ sky130_fd_sc_hd__nand2_1
X_4445_ _0786_ _0603_ _0787_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__o21ai_1
X_4376_ _3177_ _0348_ _0717_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__a211oi_1
X_7164_ _0114_ _0275_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_6115_ _0894_ _0520_ _1039_ _0524_ _2444_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__a221oi_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _0045_ _0206_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _0827_ _3407_ _0976_ _3410_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__o22ai_1
X_6948_ _3054_ _3055_ clknet_1_0__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__o21ai_2
X_6879_ _3036_ _3037_ clknet_1_0__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4230_ _3251_ _0553_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__and2_1
X_4161_ _0500_ _0504_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ _0434_ _0435_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__nand2_1
X_6802_ _2993_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4994_ _0538_ _0521_ _0442_ _0525_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__a221oi_1
X_6733_ _2925_ _2928_ vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__nand2_1
X_3945_ _3482_ vssd1 vssd1 vccd1 vccd1 _3483_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6664_ _2860_ _2861_ _2820_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__nand3_1
X_3876_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _3414_ sky130_fd_sc_hd__buf_2
X_5615_ _0488_ _0534_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6595_ _2790_ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__nand2_1
X_5546_ _0786_ _3349_ _1879_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__o21ai_1
X_5477_ _1018_ _0409_ _1809_ _1810_ _1811_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__o2111a_1
X_4428_ _0522_ _0521_ _0768_ _0525_ _0770_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__a221oi_1
X_7147_ _0097_ _0258_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
X_4359_ _3496_ _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__nand2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7078_ _0028_ _0189_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[106\]
+ sky130_fd_sc_hd__dfxtp_1
X_6029_ _0676_ _3313_ _0837_ _3317_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__3041_ clknet_0__3041_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3041_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3730_ _3267_ _3219_ vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3592_ _3142_ net32 vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__nand2_1
X_6380_ _2635_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__clkbuf_1
X_5400_ _1673_ _1734_ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__nand3_1
X_5331_ _0323_ _3296_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__nand2_1
X_5262_ _1597_ _1598_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__nand2_1
X_7001_ _3066_ _3067_ clknet_1_1__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4213_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__clkbuf_4
X_5193_ _3372_ _3452_ _3358_ _3456_ _1529_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__a221oi_1
X_4144_ _0487_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _0417_ _0418_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__nand2_1
X_6716_ _2908_ _2911_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__nand2_1
X_4977_ _0739_ _0445_ _0447_ _0435_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__a221oi_1
X_3928_ _3449_ _3452_ _3453_ _3456_ _3465_ vssd1 vssd1 vccd1 vccd1 _3466_ sky130_fd_sc_hd__a221oi_1
X_6647_ _2810_ _2844_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__nand2_1
X_3859_ _3120_ _3396_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _3397_
+ sky130_fd_sc_hd__and3_2
X_6578_ _2777_ _2752_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] egd_top.BitStream_buffer.BitStream_buffer_output\[6\]
+ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__a211o_1
X_5529_ _3244_ _3250_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4900_ _1237_ _3291_ _1238_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5880_ _0587_ _0765_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__nand2_1
X_4831_ _0412_ _3152_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nand2_1
X_4762_ _1100_ _3291_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6501_ _2714_ _2689_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__and2_1
X_3713_ _3215_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__and3_4
X_4693_ _0417_ _3163_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6432_ _2671_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
X_3644_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3575_ _3132_ _3124_ _3125_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__and3_1
X_6363_ net39 vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5314_ _3445_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _1650_
+ sky130_fd_sc_hd__nand2_1
X_6294_ _2576_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _1580_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5176_ _3386_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _1513_
+ sky130_fd_sc_hd__nand2_1
X_4127_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__buf_2
X_4058_ _3186_ _0390_ _3189_ _0393_ _0401_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _3295_ _0801_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__nand2_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6981_ _3060_ _3061_ clknet_1_0__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__o21ai_2
X_5932_ _3458_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _2263_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5863_ _0498_ _0538_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5794_ _3370_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _2126_
+ sky130_fd_sc_hd__nand2_1
X_4814_ _1150_ _1151_ _1152_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__and4_1
X_4745_ _1068_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4676_ _0967_ _0984_ _0999_ _1016_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__and4_1
X_6415_ _2659_ _2645_ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3627_ _3176_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__clkbuf_1
X_3558_ _3115_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__nand2_2
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[5] sky130_fd_sc_hd__buf_12
X_6346_ _2611_ _2601_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__and2_1
X_6277_ net16 _3395_ _2551_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__mux2_1
X_5228_ _0434_ _0731_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__nand2_1
X_5159_ _3295_ _3300_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4530_ _0817_ _0835_ _0852_ _0871_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__and4_1
X_4461_ _3245_ _3213_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7180_ _0130_ _0291_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ sky130_fd_sc_hd__dfxtp_2
X_6200_ _2511_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6131_ _0765_ _0613_ _0916_ _0617_ _2460_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__a221oi_1
X_4392_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _0649_ _3471_ _2389_ _2390_ _2391_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__o2111a_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5013_ _0577_ _0614_ _0781_ _0618_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__a221oi_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6964_ _3057_ _3058_ clknet_1_1__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__o21ai_2
X_6895_ clknet_1_0__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__buf_1
X_5915_ _0607_ _3342_ _0593_ _3346_ _2245_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__a221oi_1
X_5846_ _0394_ _0408_ _2175_ _2176_ _2177_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_90_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5777_ _0683_ _3222_ _0844_ _3228_ _2108_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__a221oi_1
X_4728_ _0563_ _0776_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4659_ _3475_ _0329_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6329_ net15 _0662_ _2470_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _3488_ _3490_ _3491_ _3493_ _3498_ vssd1 vssd1 vccd1 vccd1 _3499_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5700_ _2031_ _2032_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6680_ _2797_ _2809_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1
+ vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__o21ai_1
X_3892_ _3422_ _3424_ _3429_ vssd1 vssd1 vccd1 vccd1 _3430_ sky130_fd_sc_hd__o21ai_1
X_5631_ _1963_ _1964_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__nand2_1
X_5562_ _1518_ _3441_ _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__o21ai_1
X_4513_ _0329_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__inv_2
X_5493_ _0772_ _0486_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__o21ai_1
X_4444_ _0606_ _0593_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4375_ _0354_ egd_top.BitStream_buffer.BS_buffer\[119\] _0356_ egd_top.BitStream_buffer.BS_buffer\[120\]
+ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__a22o_1
X_7163_ _0113_ _0274_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6114_ _0743_ _0527_ _0425_ _0530_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__o22ai_1
X_7094_ _0044_ _0205_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _2364_ _2367_ _2370_ _2374_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__and4_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6947_ clknet_1_1__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__buf_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6878_ _3036_ _3037_ clknet_1_0__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__o21ai_2
X_5829_ _2150_ _2152_ _2155_ _2160_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4160_ _0503_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _0504_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4091_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__buf_2
X_6801_ _2756_ _2833_ _2760_ vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4993_ _0545_ _0528_ _0772_ _0531_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__o22ai_1
X_6732_ _2897_ _2927_ _2901_ vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__nand3_1
X_3944_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _3482_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3875_ _3395_ _3401_ _3402_ _3405_ _3412_ vssd1 vssd1 vccd1 vccd1 _3413_ sky130_fd_sc_hd__a221oi_1
X_6663_ _3111_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5614_ _1930_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__nand2_1
X_6594_ _2792_ vssd1 vssd1 vccd1 vccd1 _2793_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5545_ _3352_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _1879_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5476_ _0716_ _0422_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__or2_1
X_4427_ _0529_ _0528_ _0769_ _0531_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__o22ai_1
X_7146_ _0096_ _0257_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__clkbuf_4
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7077_ _0027_ _0188_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_4289_ _0632_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__buf_2
X_6028_ _3250_ _3280_ _3285_ _3255_ _2357_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3660_ _3201_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3591_ _3139_ _3146_ _3142_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5330_ _1664_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5261_ _0588_ _1210_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7000_ _3066_ _3067_ clknet_1_1__leaf__3068_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__o21ai_2
X_4212_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__buf_2
X_5192_ _1527_ _1528_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ _3242_ _0483_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__and2_1
X_4074_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6715_ _2909_ _2910_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__nand2_1
X_4976_ _1313_ _1314_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__nand2_1
X_3927_ _3460_ _3464_ vssd1 vssd1 vccd1 vccd1 _3465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6646_ _2842_ _2843_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3858_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _3396_ sky130_fd_sc_hd__inv_2
X_6577_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] egd_top.BitStream_buffer.BitStream_buffer_output\[2\]
+ _2750_ vssd1 vssd1 vccd1 vccd1 _2777_ sky130_fd_sc_hd__o21a_1
X_3789_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__clkbuf_4
X_5528_ _3236_ _3255_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5459_ _1790_ _1791_ _1792_ _1793_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__and4_1
X_7129_ _0079_ _0240_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4830_ _1160_ _1164_ _1166_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__and4_1
X_4761_ _3295_ _3224_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3712_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__clkbuf_4
X_6500_ net4 _1210_ _2707_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4692_ _0412_ _0733_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6431_ _2670_ _2668_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__and2_1
X_3643_ _3188_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__clkbuf_1
X_6362_ net6 _0607_ _2620_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3574_ net42 vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__inv_2
X_5313_ _3340_ _3417_ _3344_ _3421_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__a221oi_1
X_6293_ _2575_ _2559_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__and2_1
X_5244_ _0503_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _1581_
+ sky130_fd_sc_hd__nand2_1
X_5175_ _0972_ _3361_ _3376_ _3365_ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__a221oi_1
X_4126_ _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4057_ _0394_ _0396_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4959_ _3491_ _0382_ _3488_ _0385_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6629_ _2797_ _2809_ _2750_ vssd1 vssd1 vccd1 vccd1 _2827_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6980_ _3060_ _3061_ clknet_1_0__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__o21ai_2
X_5931_ _3418_ _3434_ _3437_ _3428_ _2261_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5862_ _1202_ _0485_ _2193_ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5793_ _0818_ _3342_ _0607_ _3346_ _2124_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__a221oi_1
X_4813_ _0338_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _1153_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4744_ _1072_ _1077_ _1081_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4675_ _1004_ _1006_ _1010_ _1015_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__and4_1
X_6414_ net6 _0448_ _2656_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__mux2_1
X_3626_ _3175_ _3166_ vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__and2_1
X_3557_ _3114_ vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__inv_2
X_6345_ net10 _3322_ _2469_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__mux2_1
X_6276_ _2564_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
X_5227_ _0430_ _0465_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__nand2_1
X_5158_ _1130_ _3254_ _3395_ _3258_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__a221oi_1
X_4109_ _0451_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__nand2_1
X_5089_ _3488_ _0382_ _0700_ _0385_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _3237_ _3224_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4391_ _0417_ _0733_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__nand2_1
X_6130_ _0757_ _0620_ _0908_ _0623_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_1_0__f__3065_ clknet_0__3065_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3065_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _0960_ _3484_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__or2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _1219_ _0621_ _1350_ _0624_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__o22ai_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6963_ _3057_ _3058_ clknet_1_1__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6894_ _3027_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__buf_4
X_5914_ _1215_ _3349_ _2244_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__o21ai_1
X_5845_ _1157_ _0421_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5776_ _2106_ _2107_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4727_ _1062_ _1064_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__and3_1
X_4658_ _0987_ _0990_ _0994_ _0998_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3609_ _3162_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__clkbuf_1
X_4589_ _0776_ _0556_ _0927_ _0560_ _0930_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__a221oi_1
X_6328_ _2599_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
X_6259_ _2552_ _2536_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ _3496_ _3497_ vssd1 vssd1 vccd1 vccd1 _3498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3891_ _3427_ _3428_ vssd1 vssd1 vccd1 vccd1 _3429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _0567_ _0573_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5561_ _3444_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _1895_
+ sky130_fd_sc_hd__nand2_1
X_4512_ _3480_ _3476_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5492_ _0489_ _0919_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4443_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4374_ _0716_ _0351_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nor2_1
X_7162_ _0112_ _0273_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_6113_ _2436_ _2440_ _2441_ _2442_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__and4b_1
X_7093_ _0043_ _0204_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ egd_top.BitStream_buffer.BS_buffer\[72\] _3378_ _0927_ _3382_ _2373_ vssd1
+ vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__a221oi_2
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6946_ _3027_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6877_ _3036_ _3037_ clknet_1_0__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__o21ai_2
X_5828_ _2156_ _2157_ _2158_ _2159_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__and4_1
X_5759_ _0916_ _0575_ _0518_ _0579_ _2091_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4090_ _0433_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__clkbuf_4
X_6800_ _2943_ _2991_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__nand2_1
X_4992_ _1324_ _1328_ _1329_ _1330_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__and4b_1
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6731_ _2926_ _2861_ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _3480_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _3481_
+ sky130_fd_sc_hd__nand2_1
X_3874_ _3406_ _3408_ _3409_ _3411_ vssd1 vssd1 vccd1 vccd1 _3412_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6662_ _2838_ _2859_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__nand2_1
X_5613_ _1934_ _1938_ _1942_ _1946_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6593_ _2791_ _2780_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5544_ _0551_ _3325_ _0557_ _3329_ _1877_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__a221oi_1
X_5475_ _0417_ _3183_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4426_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__inv_2
X_7145_ _0095_ _0256_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__inv_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7076_ _0026_ _0187_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[108\]
+ sky130_fd_sc_hd__dfxtp_2
X_4288_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__clkbuf_2
X_6027_ _1499_ _3290_ _2356_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__o21ai_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6929_ _3048_ _3049_ clknet_1_1__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3590_ net32 _3130_ _3127_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5260_ _0583_ _1055_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4211_ _0554_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__clkbuf_2
X_5191_ _3463_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _1528_
+ sky130_fd_sc_hd__nand2_1
X_4142_ _0485_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__clkbuf_4
X_4073_ _0416_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__buf_2
X_4975_ _0456_ egd_top.BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _1314_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _3463_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _3464_
+ sky130_fd_sc_hd__nand2_1
X_6714_ _2814_ _2750_ vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__nand2_1
X_3857_ egd_top.BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _3395_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6645_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6576_ _2776_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ sky130_fd_sc_hd__inv_2
X_3788_ _3325_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5527_ _3150_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__o21ai_1
X_5458_ _0338_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _1793_
+ sky130_fd_sc_hd__nand2_1
X_5389_ _0510_ _0576_ _0515_ _0580_ _1724_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__a221oi_1
X_4409_ _0475_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0752_
+ sky130_fd_sc_hd__nand2_1
X_7128_ _0078_ _0239_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7059_ _0009_ _0170_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4760_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3711_ _3213_ _3223_ _3224_ _3229_ _3248_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__a221oi_1
X_4691_ _1021_ _1025_ _1028_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6430_ net16 _0435_ _2656_ vssd1 vssd1 vccd1 vccd1 _2670_ sky130_fd_sc_hd__mux2_1
X_3642_ _3187_ _3166_ vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__and2_1
X_6361_ _2622_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3573_ _3127_ _3128_ _3130_ vssd1 vssd1 vccd1 vccd1 _3131_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5312_ _3348_ _3424_ _1647_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6292_ net11 _3453_ _2550_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5243_ _0499_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _1580_
+ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__3041_ _3041_ vssd1 vssd1 vccd1 vccd1 clknet_0__3041_ sky130_fd_sc_hd__clkbuf_16
X_5174_ _3348_ _3368_ _1510_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__o21ai_1
X_4125_ _3316_ _0406_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__and2_1
X_4056_ _0399_ _3192_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4958_ _3183_ _0361_ _3186_ _0364_ _1296_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a221oi_1
X_3909_ _3440_ _3442_ _3446_ vssd1 vssd1 vccd1 vccd1 _3447_ sky130_fd_sc_hd__o21ai_1
X_4889_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] _3081_ vssd1
+ vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6628_ _2745_ _2820_ _2742_ _2825_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6559_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] vssd1 vssd1 vccd1 vccd1
+ _2760_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5930_ _3422_ _3441_ _2260_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5861_ _0488_ _0442_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4812_ _0333_ _3509_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__nand2_1
X_5792_ _1078_ _3349_ _2123_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4743_ _0584_ _0614_ _0573_ _0618_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6413_ _2658_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
X_4674_ _1011_ _1012_ _1013_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__and4_1
X_3625_ net3 _3174_ _3159_ vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3556_ _3112_ _3113_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__nand2_2
X_6344_ _2610_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
X_6275_ _2563_ _2559_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5226_ _0716_ _0409_ _1560_ _1561_ _1562_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5157_ _1492_ _1493_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__nand2_1
X_4108_ egd_top.BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__clkbuf_4
X_5088_ _3186_ _0361_ _3189_ _0364_ _1425_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__a221oi_1
X_4039_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4390_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _3479_ _0648_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__nand2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__inv_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6962_ _3057_ _3058_ clknet_1_0__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__o21ai_2
X_6893_ _3024_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__buf_4
X_5913_ _3352_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _2244_
+ sky130_fd_sc_hd__nand2_1
X_5844_ _0416_ _3192_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5775_ _3244_ _3432_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__nand2_1
X_4726_ _0448_ _0537_ _0457_ _0541_ _1066_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__a221oi_1
X_4657_ _3418_ _3452_ _3428_ _3456_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__a221oi_1
X_3608_ _3160_ _3161_ vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4588_ _0928_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__nand2_1
X_6327_ _2598_ _2580_ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__and2_1
X_3539_ _3093_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__inv_2
X_6258_ net7 _3432_ _2551_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__mux2_1
X_5209_ _1535_ _1537_ _1540_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__and4_1
X_6189_ net11 _0324_ _2479_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3890_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _3428_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5560_ _3354_ _3416_ _0662_ _3420_ _1893_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__a221oi_1
X_4511_ _3475_ _0339_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__nand2_1
X_5491_ _1808_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__nand2_1
X_4442_ _0577_ _0576_ _0781_ _0580_ _0784_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__a221oi_2
X_4373_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__inv_2
X_7161_ _0111_ _0272_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_6112_ _0513_ _0739_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__nand2_1
X_7092_ _0042_ _0203_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3047_ clknet_0__3047_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3047_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _2371_ _2372_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__nand2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6945_ _3024_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6876_ _3036_ _3037_ clknet_1_0__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5827_ _0337_ egd_top.BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _2159_
+ sky130_fd_sc_hd__nand2_1
X_5758_ _2089_ _2090_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__nand2_1
X_4709_ _0731_ _0464_ _0418_ _0468_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__a221oi_1
X_5689_ _2020_ _2021_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6730_ _2913_ _2923_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__nand2_1
X_4991_ _0514_ _0768_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__nand2_1
X_3942_ _3479_ vssd1 vssd1 vccd1 vccd1 _3480_ sky130_fd_sc_hd__buf_2
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6661_ _2846_ _2858_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__nor2_1
X_3873_ _3410_ vssd1 vssd1 vccd1 vccd1 _3411_ sky130_fd_sc_hd__buf_2
X_6592_ _2781_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__inv_2
X_5612_ _3174_ _0463_ _3177_ _0467_ _1945_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5543_ _0622_ _3122_ _1876_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5474_ _0412_ _3177_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__nand2_1
X_4425_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__buf_2
XFILLER_0_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7144_ _0094_ _0255_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_4356_ _0693_ _3472_ _0694_ _0696_ _0698_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__o2111a_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _0025_ _0186_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[109\]
+ sky130_fd_sc_hd__dfxtp_1
X_4287_ _0630_ _3120_ _3396_ _3218_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__and4b_1
X_6026_ _3294_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _2356_
+ sky130_fd_sc_hd__nand2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6928_ _3048_ _3049_ clknet_1_1__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6859_ _3033_ _3034_ clknet_1_0__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4210_ _3217_ _0553_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__and2_1
X_5190_ _3459_ _0840_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__nand2_1
X_4141_ _3234_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__nand2_2
X_4072_ _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__clkbuf_2
X_4974_ _0451_ _0894_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nand2_1
X_6713_ _2797_ _2809_ _2754_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__o21ai_1
X_3925_ _3462_ vssd1 vssd1 vccd1 vccd1 _3463_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6644_ _2841_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3856_ _3339_ _3357_ _3375_ _3393_ vssd1 vssd1 vccd1 vccd1 _3394_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6575_ _2740_ _2745_ _2775_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3787_ _3324_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5526_ _1738_ _1860_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__nor2_1
X_5457_ _0333_ _3296_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4408_ _0471_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _0751_
+ sky130_fd_sc_hd__nand2_1
X_5388_ _1722_ _1723_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__nand2_1
X_7127_ _0077_ _0238_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_4339_ _3418_ _3417_ _3428_ _3421_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7058_ _0008_ _0169_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[87\]
+ sky130_fd_sc_hd__dfxtp_1
X_6009_ _0515_ _0613_ _0765_ _0617_ _2339_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3710_ _3239_ _3247_ vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4690_ _3195_ _0390_ _3199_ _0393_ _1030_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__a221oi_1
X_3641_ net14 _3186_ _3159_ vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3572_ _3129_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__inv_2
X_6360_ _2621_ _2601_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5311_ _3427_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _1647_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6291_ _2574_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
X_5242_ _0542_ _0486_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__o21ai_1
X_5173_ _3371_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _1510_
+ sky130_fd_sc_hd__nand2_1
X_4124_ _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__clkbuf_4
Xinput1 la_data_in_47_32[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
X_4055_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__buf_2
X_4957_ _0349_ _0367_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__o21ai_1
X_3908_ _3445_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _3446_
+ sky130_fd_sc_hd__nand2_1
X_4888_ _1091_ _1227_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6627_ _2824_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__inv_2
X_3839_ _3302_ _3323_ vssd1 vssd1 vccd1 vccd1 _3377_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6558_ _2757_ _2758_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__nand2_1
X_6489_ _3156_ net42 _2474_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__nand3_4
X_5509_ _0577_ _0556_ _0781_ _0560_ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a221oi_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5860_ _2174_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4811_ _0328_ _0865_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nand2_1
X_5791_ _3352_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _2123_
+ sky130_fd_sc_hd__nand2_1
X_4742_ _0941_ _0621_ _1082_ _0624_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4673_ _0338_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1014_
+ sky130_fd_sc_hd__nand2_1
X_6412_ _2657_ _2645_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3624_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3555_ _3111_ egd_top.BitStream_buffer.pc_previous\[0\] vssd1 vssd1 vccd1 vccd1 _3113_
+ sky130_fd_sc_hd__nand2_4
X_6343_ _2609_ _2601_ vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__and2_1
X_6274_ net2 _1130_ _2551_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5225_ _1161_ _0422_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5156_ _3270_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _1493_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4107_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__buf_2
X_5087_ _0716_ _0367_ _1424_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__o21ai_1
X_4038_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _0508_ _0452_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _0557_ _0596_ _0776_ _0600_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__a221oi_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6961_ _3057_ _3058_ clknet_1_1__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__o21ai_2
X_6892_ _3039_ _3040_ clknet_1_0__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__o21ai_2
X_5912_ _0927_ _3325_ _0611_ _3329_ _2242_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5843_ _0411_ _3186_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5774_ _3236_ _3439_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4725_ _0923_ _0544_ _1065_ _0547_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4656_ _0995_ _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__nand2_1
X_3607_ _3080_ vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__buf_6
X_4587_ _0568_ _0551_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__nand2_1
X_3538_ _3097_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_1
X_6326_ net16 _3354_ _2470_ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6257_ _2550_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__clkbuf_4
X_5208_ _1541_ _1542_ _1543_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__and4_1
X_6188_ _2503_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__clkbuf_1
X_5139_ _0776_ _0596_ _0927_ _0600_ _1476_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4510_ _0839_ _0843_ _0847_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__and4_1
X_5490_ _1812_ _1816_ _1820_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4441_ _0782_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__nand2_1
X_7160_ _0110_ _0271_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_6111_ _0508_ _0746_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__nand2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _0656_ _0674_ _0692_ _0714_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__and4_1
X_7091_ _0041_ _0202_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _3389_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _2372_
+ sky130_fd_sc_hd__nand2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6944_ _3051_ _3052_ clknet_1_1__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6875_ _3036_ _3037_ clknet_1_0__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__o21ai_2
X_5826_ _0332_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _2158_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5757_ _0587_ _0515_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__nand2_1
X_4708_ _1047_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__nand2_1
X_5688_ _3462_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _2021_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4639_ _3386_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _0980_
+ sky130_fd_sc_hd__nand2_1
X_6309_ _2586_ _2580_ vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4990_ _0509_ _0522_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__nand2_1
X_3941_ _3478_ vssd1 vssd1 vccd1 vccd1 _3479_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6660_ _2854_ _2857_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3872_ _3234_ _3398_ vssd1 vssd1 vccd1 vccd1 _3410_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6591_ _2779_ _2789_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5611_ _1943_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__nand2_1
X_5542_ _3334_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _1876_
+ sky130_fd_sc_hd__nand2_1
X_5473_ _1799_ _1802_ _1804_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__and4_1
X_4424_ _0759_ _0763_ _0764_ _0766_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__and4b_1
X_7143_ _0093_ _0254_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_4355_ _0697_ _3485_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__or2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7074_ _0024_ _0185_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4286_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] egd_top.BitStream_buffer.pc\[1\]
+ _3115_ _3470_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__o41a_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _3414_ _3253_ _3418_ _3257_ _2354_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__a221oi_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6927_ _3048_ _3049_ clknet_1_0__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6858_ _3033_ _3034_ clknet_1_0__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5809_ _3414_ _3434_ _3437_ _3418_ _2140_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__a221oi_1
X_6789_ _2965_ _2981_ _2967_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4140_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__clkbuf_4
X_4071_ _3251_ _0407_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _1308_ _0427_ _1309_ _1310_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__o2111a_1
X_6712_ _2875_ _2817_ _2831_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__nand3_1
X_3924_ _3461_ vssd1 vssd1 vccd1 vccd1 _3462_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6643_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3855_ _3376_ _3379_ _3380_ _3383_ _3392_ vssd1 vssd1 vccd1 vccd1 _3393_ sky130_fd_sc_hd__a221oi_1
X_6574_ _2773_ _2774_ vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__nand2_1
X_3786_ _3267_ _3323_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__and2_1
X_5525_ _3212_ _1859_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ _0328_ _0648_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4407_ _0448_ _0445_ _0447_ _0457_ _0749_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__a221oi_1
X_5387_ _0588_ _1055_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__nand2_1
X_7126_ _0076_ _0237_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_4338_ _3366_ _3424_ _0680_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__o21ai_1
X_7057_ _0007_ _0168_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[88\]
+ sky130_fd_sc_hd__dfxtp_1
X_4269_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__clkbuf_2
X_6008_ _0481_ _0620_ _0757_ _0623_ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3640_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__buf_2
X_3571_ _3103_ _3107_ vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__nor2_1
X_6290_ _2573_ _2559_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__and2_1
X_5310_ _3428_ _3401_ _0679_ _3405_ _1645_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5241_ _0489_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _1578_
+ sky130_fd_sc_hd__nand2_1
X_5172_ _3380_ _3343_ _3322_ _3347_ _1508_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__a221oi_1
X_4123_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__clkbuf_2
X_4054_ _0397_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__clkbuf_2
Xinput2 la_data_in_47_32[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_4
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4956_ _0370_ _3180_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__nand2_1
X_3907_ _3444_ vssd1 vssd1 vccd1 vccd1 _3445_ sky130_fd_sc_hd__buf_2
X_4887_ _3212_ _1226_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6626_ _2740_ _2822_ _2823_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__or3_1
X_3838_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _3376_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6557_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] vssd1 vssd1 vccd1 vccd1
+ _2758_ sky130_fd_sc_hd__inv_2
X_3769_ _3301_ _3116_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__nor2_4
X_5508_ _1841_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__nand2_1
X_6488_ _3090_ _3114_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__nor2_1
X_5439_ _1391_ _3442_ _1773_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__o21ai_1
X_7109_ _0059_ _0220_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4810_ _0323_ _3512_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5790_ _0776_ _3325_ _0927_ _3329_ _2121_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4741_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4672_ _0333_ _0865_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nand2_1
X_6411_ net7 _0442_ _2656_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__mux2_1
X_3623_ _3173_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ egd_top.BitStream_buffer.pc_previous\[0\] _3111_ vssd1 vssd1 vccd1 vccd1 _3112_
+ sky130_fd_sc_hd__or2_1
X_6342_ net11 _3380_ _2469_ vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__mux2_1
X_6273_ _2562_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5224_ _0417_ _3177_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__nand2_1
X_5155_ _3263_ _0991_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4106_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__clkbuf_2
X_5086_ _0370_ _3183_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4037_ _3267_ _0345_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _0919_ _0493_ _0495_ _0534_ _2318_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4939_ _1002_ _3472_ _1275_ _1276_ _1277_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__o2111a_1
XANTENNA_40 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6609_ _2793_ _2798_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__3062_ clknet_0__3062_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3062_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6960_ clknet_1_1__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__buf_1
X_5911_ _1082_ _3122_ _2241_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6891_ _3039_ _3040_ clknet_1_0__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5842_ _2165_ _2168_ _2170_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5773_ _3150_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__inv_2
X_4655_ _3463_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _0996_
+ sky130_fd_sc_hd__nand2_1
X_3606_ net7 _3152_ _3159_ vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__mux2_1
X_4586_ _0563_ _0557_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3537_ _3095_ _3080_ _3096_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__and3_1
X_6325_ _2597_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6256_ _2471_ _3132_ _2475_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__nand3_4
X_5207_ _0338_ _3512_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nand2_1
X_6187_ _2502_ _2492_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__and2_1
X_5138_ _1474_ _0603_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__o21ai_1
X_5069_ _3503_ _3485_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4440_ _0588_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _0783_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6110_ _0534_ _0493_ _0495_ _0538_ _2439_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__a221oi_1
X_4371_ _0699_ _0703_ _0707_ _0713_ vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__and4_1
X_7090_ _0040_ _0201_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _3385_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _2371_
+ sky130_fd_sc_hd__nand2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6943_ _3051_ _3052_ clknet_1_1__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__o21ai_2
X_6874_ _3036_ _3037_ clknet_1_0__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5825_ _0327_ _3238_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5756_ _0582_ _0765_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4707_ _0475_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _1048_
+ sky130_fd_sc_hd__nand2_1
X_5687_ _3458_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _2020_
+ sky130_fd_sc_hd__nand2_1
X_4638_ _3344_ _3361_ _3354_ _3365_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ _0499_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0911_
+ sky130_fd_sc_hd__nand2_1
X_6308_ net7 _0840_ _2470_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__mux2_1
X_6239_ _2538_ _2536_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__and2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ _3242_ _3469_ vssd1 vssd1 vccd1 vccd1 _3478_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3871_ egd_top.BitStream_buffer.BS_buffer\[37\] vssd1 vssd1 vccd1 vccd1 _3409_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6590_ _2788_ _2750_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__nand2_1
X_5610_ _0474_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _1944_
+ sky130_fd_sc_hd__nand2_1
X_5541_ _1865_ _1869_ _1872_ _1874_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5472_ _0796_ _0390_ _0947_ _0393_ _1806_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__a221oi_1
X_4423_ _0514_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__nand2_1
X_7142_ _0092_ _0253_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_4354_ _0339_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__inv_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7073_ _0023_ _0184_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[111\]
+ sky130_fd_sc_hd__dfxtp_1
X_6024_ _2352_ _2353_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__nand2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _0480_ _0628_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__nor2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6926_ _3048_ _3049_ clknet_1_1__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6857_ _3033_ _3034_ clknet_1_0__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__o21ai_2
X_6788_ _2979_ vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__inv_2
X_5808_ _1767_ _3441_ _2139_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__o21ai_1
X_5739_ _1065_ _0485_ _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4070_ _0412_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nand2_1
X_4972_ _1037_ _0439_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__or2_1
X_6711_ _2903_ _2875_ _2906_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__nand3_1
X_3923_ _3312_ _3397_ vssd1 vssd1 vccd1 vccd1 _3461_ sky130_fd_sc_hd__and2_1
X_6642_ _2807_ _2839_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3854_ _3387_ _3391_ vssd1 vssd1 vccd1 vccd1 _3392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6573_ _3149_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] vssd1 vssd1
+ vccd1 vccd1 _2774_ sky130_fd_sc_hd__nor2_1
X_3785_ _3121_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__buf_2
X_5524_ _1796_ _1857_ _1858_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__nand3_2
X_5455_ _0323_ _3246_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4406_ _0747_ _0748_ vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nand2_1
X_7125_ _0075_ _0236_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_5386_ _0583_ _1192_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _3427_ _0679_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__nand2_1
X_7056_ _0006_ _0167_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[89\]
+ sky130_fd_sc_hd__dfxtp_1
X_4268_ _3302_ _0552_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__and2_1
X_6007_ _0577_ _0595_ _0781_ _0599_ _2337_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__a221oi_1
X_4199_ _3267_ _0484_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__nand2_2
XFILLER_0_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6909_ _3045_ _3046_ clknet_1_0__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3570_ _3101_ net33 net32 vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__or3b_1
XFILLER_0_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _1559_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5171_ _1506_ _3350_ _1507_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__o21ai_1
X_4122_ _3307_ _0407_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__and2_1
X_4053_ _3302_ _0344_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__and2_1
Xinput3 la_data_in_47_32[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_4
X_4955_ _3189_ _0348_ _1292_ _1293_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3906_ _3443_ vssd1 vssd1 vccd1 vccd1 _3444_ sky130_fd_sc_hd__clkbuf_2
X_4886_ _1156_ _1224_ _1225_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__nand3_2
X_6625_ _2775_ _2784_ _2794_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__and3_1
X_3837_ _3358_ _3361_ _3362_ _3365_ _3374_ vssd1 vssd1 vccd1 vccd1 _3375_ sky130_fd_sc_hd__a221oi_1
X_3768_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__clkbuf_4
X_6556_ _2755_ _2756_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__nand2_1
X_5507_ _0568_ _0584_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__nand2_1
X_3699_ _3236_ vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__buf_2
X_6487_ _3230_ _3090_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5438_ _3445_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _1773_
+ sky130_fd_sc_hd__nand2_1
X_5369_ _0545_ _0486_ _1704_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__o21ai_1
X_7108_ _0058_ _0219_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_7039_ _3075_ _3076_ clknet_1_1__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__o21ai_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4740_ _0564_ _0596_ _0551_ _0600_ _1080_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_83_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4671_ _0328_ _0708_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6410_ _2655_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__clkbuf_4
X_3622_ _3172_ _3166_ vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6341_ _2608_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__clkbuf_1
X_3553_ _3109_ _3110_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__nand2_2
X_6272_ _2561_ _2559_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__and2_1
X_5223_ _0412_ _3171_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__nand2_1
X_5154_ _3264_ _3223_ _3250_ _3229_ _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__a221oi_1
X_4105_ _3292_ _0406_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__and2_1
X_5085_ _3192_ _0348_ _1421_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4036_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _2316_ _2317_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4938_ _3500_ _3485_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4869_ _0611_ _0556_ _0615_ _0560_ _1208_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a221oi_1
XANTENNA_41 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_30 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6608_ _2799_ _2752_ _2805_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__a21oi_1
X_6539_ _3111_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ _3334_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _2241_
+ sky130_fd_sc_hd__nand2_1
X_6890_ _3039_ _3040_ clknet_1_1__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5841_ _0701_ _0389_ _0695_ _0392_ _2172_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5772_ _1983_ _2104_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4723_ _0919_ _0521_ _0534_ _0525_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4654_ _3459_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _0995_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4585_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__clkbuf_4
X_3605_ _3158_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__clkbuf_4
X_3536_ _3094_ net36 vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__nand2_1
X_6324_ _2596_ _2580_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__and2_1
X_6255_ _2549_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5206_ _0333_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _1543_
+ sky130_fd_sc_hd__nand2_1
X_6186_ net12 _0334_ _2479_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__mux2_1
X_5137_ _0606_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _1475_
+ sky130_fd_sc_hd__nand2_1
X_5068_ _3480_ _0334_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__nand2_1
X_4019_ _0362_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4370_ _0709_ _0710_ _0711_ _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__and4_1
Xclkbuf_1_0__f__3044_ clknet_0__3044_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3044_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _0818_ _3360_ _0607_ _3364_ _2369_ vssd1 vssd1 vccd1 vccd1 _2370_ sky130_fd_sc_hd__a221oi_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ _3051_ _3052_ clknet_1_1__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6873_ _3036_ _3037_ clknet_1_1__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5824_ _0322_ _3224_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5755_ _0932_ _0555_ _1073_ _0559_ _2087_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__a221oi_1
X_4706_ _0471_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1047_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5686_ _3453_ _3434_ _3437_ _3414_ _2018_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4637_ _0976_ _3368_ _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4568_ _0908_ _0486_ _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__o21ai_1
X_3519_ _3080_ vssd1 vssd1 vccd1 vccd1 _3081_ sky130_fd_sc_hd__buf_2
X_4499_ _3427_ _0840_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__nand2_1
X_6307_ _2585_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
X_6238_ net12 _3300_ _2515_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__mux2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _2490_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__clkbuf_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3870_ _3407_ vssd1 vssd1 vccd1 vccd1 _3408_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5540_ _0991_ _3304_ _1130_ _3309_ _1873_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5471_ _0858_ _0396_ _1805_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o21ai_1
X_4422_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__buf_2
X_7210_ _0160_ _0321_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7141_ _0091_ _0252_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4353_ _3480_ _0695_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__nand2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _0550_ _0627_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__nand2_1
X_7072_ _0022_ _0183_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_6023_ _3269_ _3449_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__nand2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6925_ _3048_ _3049_ clknet_1_0__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6856_ clknet_1_0__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__buf_1
XFILLER_0_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6787_ _2968_ _2979_ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3999_ _3321_ _3394_ _3467_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__and4_1
X_5807_ _3444_ _0679_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__nand2_1
X_5738_ _0488_ _0538_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5669_ _0937_ _3349_ _2001_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4971_ _0434_ _0465_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__nand2_1
X_3922_ _3459_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _3460_
+ sky130_fd_sc_hd__nand2_1
X_6710_ _2904_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__nand2_1
X_6641_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__xnor2_1
X_3853_ _3390_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _3391_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6572_ _2771_ _2772_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__nand2_2
X_3784_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5523_ _0633_ _0329_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__nand2_1
X_5454_ _1787_ _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__nor2_1
X_4405_ _0456_ egd_top.BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _0748_
+ sky130_fd_sc_hd__nand2_1
X_5385_ _0573_ _0556_ _0577_ _0560_ _1720_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__a221oi_1
X_7124_ _0074_ _0235_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_4336_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__buf_2
X_7055_ _0005_ _0166_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[90\]
+ sky130_fd_sc_hd__dfxtp_1
X_4267_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__clkbuf_4
X_4198_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__inv_2
X_6006_ _1219_ _0602_ _2336_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6908_ clknet_1_1__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__buf_1
XFILLER_0_49_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6839_ _3027_ vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5170_ _3353_ _3327_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__nand2_1
X_4121_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__buf_2
X_4052_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__buf_2
Xinput4 la_data_in_47_32[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_4
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4954_ _0354_ egd_top.BitStream_buffer.BS_buffer\[123\] _0356_ _3199_ vssd1 vssd1
+ vccd1 vccd1 _1293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3905_ _3292_ _3397_ vssd1 vssd1 vccd1 vccd1 _3443_ sky130_fd_sc_hd__and2_1
X_4885_ _0633_ _0701_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6624_ _2781_ _2821_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _3366_ _3368_ _3373_ vssd1 vssd1 vccd1 vccd1 _3374_ sky130_fd_sc_hd__o21ai_1
X_3767_ _3304_ vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6555_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] vssd1 vssd1 vccd1 vccd1
+ _2756_ sky130_fd_sc_hd__inv_2
X_5506_ _0563_ _0573_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3698_ _3235_ vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__clkbuf_2
X_6486_ _3113_ _2705_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[1\] sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5437_ _3344_ _3417_ _3354_ _3421_ _1771_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5368_ _0489_ _0768_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7107_ _0057_ _0218_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_5299_ _3322_ _3343_ _3327_ _3347_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__a221oi_1
X_4319_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__buf_2
X_7038_ clknet_1_0__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__buf_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4670_ _0323_ _3509_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__nand2_1
X_3621_ net4 _3171_ _3159_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__mux2_1
X_3552_ net17 vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__inv_2
X_6340_ _2607_ _2601_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6271_ net3 _0991_ _2551_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5222_ _1550_ _1553_ _1555_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__and4_1
X_5153_ _1488_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__nand2_1
X_4104_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _0354_ egd_top.BitStream_buffer.BS_buffer\[124\] _0356_ _3202_ vssd1 vssd1
+ vccd1 vccd1 _1422_ sky130_fd_sc_hd__a22o_1
X_4035_ _0378_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _0502_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _2317_
+ sky130_fd_sc_hd__nand2_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4937_ _3480_ _0329_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_31 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _1206_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__nand2_1
XANTENNA_20 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6607_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] _2801_ _2804_ vssd1
+ vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__o21ai_1
XANTENNA_42 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3819_ _3340_ _3343_ _3344_ _3347_ _3356_ vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__a221oi_1
X_4799_ _3475_ _0334_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6538_ _2739_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_6469_ _2696_ _2697_ _2698_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5840_ _3483_ _0395_ _2171_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5771_ _3149_ _2103_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__nor2_1
X_4722_ _0920_ _0528_ _0542_ _0531_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4653_ _0844_ _3435_ _3438_ _0991_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__a221oi_1
X_4584_ _0918_ _0922_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__and3_1
X_3604_ _3157_ vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3535_ net36 _3094_ vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__or2_1
X_6323_ net2 _3344_ _2470_ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__mux2_1
X_6254_ _2548_ _2536_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5205_ _0328_ _3275_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6185_ _2501_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__clkbuf_1
X_5136_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__inv_2
X_5067_ _3475_ _0708_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__nand2_1
X_4018_ _3292_ _0345_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5969_ _0429_ _3163_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6941_ _3051_ _3052_ clknet_1_1__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6872_ _3036_ _3037_ clknet_1_1__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5823_ _2153_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5754_ _2085_ _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__nand2_1
X_4705_ _0452_ _0445_ _0447_ _0746_ _1045_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__a221oi_1
X_5685_ _1644_ _3441_ _2017_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4636_ _3371_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _0977_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4567_ _0489_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0909_
+ sky130_fd_sc_hd__nand2_1
X_6306_ _2584_ _2580_ vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__and2_1
X_3518_ _3079_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__buf_6
X_4498_ egd_top.BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__buf_2
X_6237_ _2537_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _2489_ _3197_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _0509_ _0768_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__nand2_1
X_6099_ _0470_ _3183_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5470_ _0399_ _3497_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__nand2_1
X_4421_ _0509_ _0515_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7140_ _0090_ _0251_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_4352_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__clkbuf_4
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4283_ _0572_ _0592_ _0610_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__and4_1
X_7071_ _0021_ _0182_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6022_ _3262_ _3453_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__nand2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _3048_ _3049_ clknet_1_0__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6855_ _3027_ vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__buf_4
X_6786_ _2978_ _2861_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5806_ _0823_ _3416_ _0972_ _3420_ _2137_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__a221oi_1
X_3998_ _3487_ _3499_ _3514_ _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5737_ _2052_ _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__nand2_1
X_5668_ _3352_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _2001_
+ sky130_fd_sc_hd__nand2_1
X_4619_ egd_top.BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__inv_2
X_5599_ _0873_ _0421_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _0430_ _1039_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nand2_1
X_3921_ _3458_ vssd1 vssd1 vccd1 vccd1 _3459_ sky130_fd_sc_hd__buf_2
X_6640_ _2832_ _2837_ _2818_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__nand3_1
X_3852_ _3389_ vssd1 vssd1 vccd1 vccd1 _3390_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6571_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] egd_top.BitStream_buffer.BitStream_buffer_output\[14\]
+ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__nor2_1
X_3783_ _3249_ _3274_ _3299_ _3320_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5522_ _1826_ _1856_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5453_ _3508_ egd_top.BitStream_buffer.BS_buffer\[23\] _3511_ _0639_ vssd1 vssd1
+ vccd1 vccd1 _1788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4404_ _0451_ _0746_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__nand2_1
X_5384_ _1718_ _1719_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4335_ _3402_ _3401_ _0675_ _3405_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7123_ _0073_ _0234_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_7054_ _0004_ _0165_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[91\]
+ sky130_fd_sc_hd__dfxtp_1
X_4266_ _0593_ _0596_ _0597_ _0600_ _0609_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6005_ _0605_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _2336_
+ sky130_fd_sc_hd__nand2_1
X_4197_ _0540_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6907_ _3027_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6838_ _3026_ vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__buf_4
X_6769_ _2961_ _2869_ _2962_ vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3077_ clknet_0__3077_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3077_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4120_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__buf_2
X_4051_ _3307_ _0345_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__nand2_2
Xinput5 la_data_in_47_32[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4953_ _1291_ _0351_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3904_ _3441_ vssd1 vssd1 vccd1 vccd1 _3442_ sky130_fd_sc_hd__clkbuf_4
X_6623_ _2779_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__inv_2
X_4884_ _1189_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3835_ _3371_ _3372_ vssd1 vssd1 vccd1 vccd1 _3373_ sky130_fd_sc_hd__nand2_1
X_6554_ _2753_ _2754_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__nand2_1
X_3766_ _3303_ vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__clkbuf_2
X_6485_ _2704_ _2692_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__and2_1
X_5505_ _1835_ _1837_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3697_ _3234_ _3219_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__and2_1
X_5436_ _0661_ _3424_ _1770_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__o21ai_1
X_5367_ _1685_ _1702_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7106_ _0056_ _0217_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_5298_ _3331_ _3350_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__o21ai_1
X_4318_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__inv_2
X_7037_ _3026_ vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__buf_4
X_4249_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__buf_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3620_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3551_ net18 vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__inv_2
X_6270_ _2560_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5221_ _3208_ _0390_ _0634_ _0393_ _1557_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__a221oi_1
X_5152_ _3245_ _3306_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__nand2_1
X_4103_ _0446_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__clkbuf_4
X_5083_ _0394_ _0351_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__nor2_1
X_4034_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5985_ _0498_ _0442_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__nand2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4936_ _3475_ _0324_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_1
XANTENNA_32 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _0568_ _0776_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__nand2_1
XANTENNA_10 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6606_ _2803_ _2763_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3818_ _3348_ _3350_ _3355_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__o21ai_1
X_6537_ _2738_ _3080_ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__and2_1
X_4798_ _1126_ _1129_ _1133_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__and4_1
X_3749_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__clkbuf_4
X_6468_ egd_top.BitStream_buffer.pc_previous\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6399_ _2648_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
X_5419_ _0619_ _3332_ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5770_ _2040_ _2101_ _2102_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__nand3_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4721_ _1054_ _1059_ _1060_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__and4b_1
XFILLER_0_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4652_ _3409_ _3442_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__o21ai_1
X_3603_ _3132_ _3124_ _3125_ _3156_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__or4b_2
XFILLER_0_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4583_ _0442_ _0537_ _0448_ _0541_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__a221oi_2
X_3534_ _3091_ _3093_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__nor2_1
X_6322_ _2595_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
X_6253_ net1 _3255_ _2515_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__mux2_1
X_5204_ _0323_ _0648_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__nand2_1
X_6184_ _2492_ _2500_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__and2_1
X_5135_ _1055_ _0576_ _1192_ _0580_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5066_ _1393_ _1396_ _1399_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__buf_2
X_5968_ _0380_ _0408_ _2296_ _2297_ _2298_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__o2111a_1
X_4919_ _1256_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__nand2_1
X_5899_ _0844_ _3222_ _0991_ _3228_ _2229_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6940_ _3051_ _3052_ clknet_1_0__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6871_ _3036_ _3037_ clknet_1_1__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__o21ai_2
X_5822_ _3507_ egd_top.BitStream_buffer.BS_buffer\[26\] _3510_ egd_top.BitStream_buffer.BS_buffer\[27\]
+ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5753_ _0567_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _2086_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4704_ _1043_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5684_ _3444_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _2017_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4566_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3517_ net20 net22 _3078_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__o21a_4
X_6305_ net1 _0679_ _2550_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__mux2_1
X_4497_ _0675_ _3401_ _0836_ _3405_ _0838_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__a221oi_1
X_6236_ _2535_ _2536_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__and2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ net3 _0701_ _2480_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _0510_ _0494_ _0496_ _0515_ _1455_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__a221oi_1
X_6098_ _0418_ _0444_ _0446_ _0733_ _2427_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__a221oi_1
X_5049_ _3390_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _1387_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4420_ egd_top.BitStream_buffer.BS_buffer\[81\] _0494_ _0496_ egd_top.BitStream_buffer.BS_buffer\[82\]
+ _0762_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4351_ _3475_ _3482_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__nand2_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _0611_ _0614_ _0615_ _0618_ _0625_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__a221oi_1
X_7070_ _0020_ _0181_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_6021_ _0991_ _3222_ _1130_ _3228_ _2350_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__a221oi_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6923_ _3048_ _3049_ clknet_1_0__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _3024_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6785_ _2975_ _2977_ vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__nand2_1
X_5805_ _1111_ _3423_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__o21ai_1
X_3997_ _0325_ _0330_ _0335_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5736_ _2056_ _2060_ _2064_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__and4_1
X_5667_ _0557_ _3325_ _0776_ _3329_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__a221oi_1
X_4618_ _3439_ _3254_ _0683_ _3258_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5598_ _0416_ _3186_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__nand2_1
X_4549_ _0720_ _0409_ _0888_ _0889_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__o2111a_1
X_6219_ net3 _3246_ _2516_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__mux2_1
X_7199_ _0149_ _0310_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3920_ _3457_ vssd1 vssd1 vccd1 vccd1 _3458_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3851_ _3388_ vssd1 vssd1 vccd1 vccd1 _3389_ sky130_fd_sc_hd__clkbuf_2
X_3782_ _3300_ _3305_ _3306_ _3310_ _3319_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__a221oi_1
X_6570_ _2769_ _2770_ vssd1 vssd1 vccd1 vccd1 _2771_ sky130_fd_sc_hd__nand2_1
X_5521_ _1840_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5452_ _0960_ _3502_ _1100_ _3505_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__o22ai_1
X_4403_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__clkbuf_4
X_5383_ _0568_ _0589_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__nand2_1
X_4334_ _3409_ _3408_ _0676_ _3411_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__o22ai_1
X_7122_ _0072_ _0233_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_7053_ _0003_ _0164_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[92\]
+ sky130_fd_sc_hd__dfxtp_1
X_6004_ _0522_ _0575_ _0768_ _0579_ _2334_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__a221oi_1
X_4265_ _0601_ _0603_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__o21ai_1
X_4196_ _0539_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6906_ _3024_ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__buf_4
X_6837_ net21 vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6768_ _2960_ _2955_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6699_ _2860_ _2895_ _2861_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5719_ _2043_ _2046_ _2048_ _2051_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4050_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
Xinput6 la_data_in_47_32[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_4
XFILLER_0_78_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4952_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4883_ _1205_ _1222_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3903_ _3289_ _3398_ vssd1 vssd1 vccd1 vccd1 _3441_ sky130_fd_sc_hd__nand2_2
X_6622_ _2806_ _2812_ _2819_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__nand3_2
X_3834_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _3372_ sky130_fd_sc_hd__buf_2
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3765_ _3302_ _3219_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__and2_1
X_6553_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1 vccd1
+ _2754_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6484_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__or2_1
X_3696_ _3233_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__clkbuf_8
X_5504_ _0741_ _0537_ _0894_ _0541_ _1838_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__a221oi_1
X_5435_ _3427_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _1770_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5366_ _1689_ _1693_ _1697_ _1701_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__and4_1
X_7105_ _0055_ _0216_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_5297_ _3353_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _1633_
+ sky130_fd_sc_hd__nand2_1
X_4317_ _3327_ _3326_ _3336_ _3330_ _0659_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__a221oi_1
X_7036_ _3023_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__buf_4
X_4248_ _0573_ _0576_ _0577_ _0580_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__a221oi_1
X_4179_ _3307_ _0484_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__and2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3550_ _3107_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__3059_ clknet_0__3059_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3059_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5220_ _3488_ _0396_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__o21ai_1
X_5151_ _3237_ _3271_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__nand2_1
X_4102_ _0405_ _3282_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__nor2_2
X_5082_ _1374_ _1390_ _1404_ _1419_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__and4_1
X_4033_ _3119_ _0345_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _1334_ _0485_ _2314_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__o21ai_1
X_4935_ _1263_ _1266_ _1269_ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_22 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _0563_ _0927_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__nand2_1
XANTENNA_44 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6605_ _2773_ _2774_ _2802_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_33 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _3353_ _3354_ vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__nand2_1
X_4797_ _3428_ _3452_ _0679_ _3456_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__a221oi_1
X_3748_ _3285_ vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__buf_2
X_6536_ net1 _0538_ _2706_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6467_ egd_top.BitStream_buffer.pc_previous\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__or2_1
X_3679_ _3215_ egd_top.BitStream_buffer.pc\[2\] _3216_ vssd1 vssd1 vccd1 vccd1 _3217_
+ sky130_fd_sc_hd__and3_4
X_6398_ _2647_ _2645_ vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__and2_1
X_5418_ _3335_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _1753_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5349_ _1676_ _1679_ _1681_ _1684_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__and4_1
X_7019_ _3069_ _3070_ clknet_1_0__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4720_ _0514_ _0518_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__nand2_1
X_4651_ _3445_ egd_top.BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _0992_
+ sky130_fd_sc_hd__nand2_1
Xinput20 la_data_in_65 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
X_3602_ _3153_ _3154_ _3098_ _3155_ vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__a22o_2
XFILLER_0_71_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4582_ _0772_ _0544_ _0923_ _0547_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3533_ _3084_ _3092_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6321_ _2594_ _2580_ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__and2_1
X_6252_ _2547_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5203_ _1538_ _1539_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6183_ net13 _0329_ _2480_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5134_ _1470_ _1471_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__nand2_1
X_5065_ _0840_ _3452_ _3372_ _3456_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4016_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__clkbuf_2
X_5967_ _1291_ _0421_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__or2_1
X_4918_ _3390_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _1257_
+ sky130_fd_sc_hd__nand2_1
X_5898_ _2227_ _2228_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4849_ _1170_ _1188_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nand2_1
X_6519_ _2726_ _3080_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__3041_ clknet_0__3041_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3041_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6870_ _3036_ _3037_ clknet_1_1__leaf__3038_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5821_ _3311_ _3501_ _3315_ _3504_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5752_ _0562_ _0781_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4703_ _0456_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _1044_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5683_ _0662_ _3416_ _0823_ _3420_ _2015_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4634_ _0662_ _3343_ _0823_ _3347_ _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4565_ _0887_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3516_ net23 net22 vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__or2b_4
X_6304_ _2583_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
X_4496_ _0676_ _3408_ _0837_ _3411_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__o22ai_1
X_6235_ _3165_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__buf_6
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _2488_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _1453_ _1454_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__nand2_1
X_6097_ _2425_ _2426_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__nand2_1
X_5048_ _3386_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _1386_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6999_ clknet_1_0__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__buf_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4350_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__inv_2
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ _0619_ _0621_ _0622_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__o22ai_1
X_6020_ _2348_ _2349_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__nand2_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6922_ _3048_ _3049_ clknet_1_0__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__o21ai_2
X_6853_ _3025_ _3028_ clknet_1_0__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__o21ai_2
X_5804_ _3426_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _2136_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6784_ _2766_ _2949_ _2976_ _2952_ vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__a211o_1
X_3996_ _0338_ _0339_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__nand2_1
X_5735_ _3177_ _0463_ _3180_ _0467_ _2067_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__a221oi_1
X_5666_ _0790_ _3122_ _1998_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__o21ai_1
X_4617_ _0956_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5597_ _0411_ _3180_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__nand2_1
X_4548_ _0404_ _0422_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__or2_1
X_4479_ _3336_ _3326_ _0657_ _3330_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__a221oi_1
X_6218_ _2524_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
X_7198_ _0148_ _0309_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _2473_ _2476_ _3089_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3850_ _3312_ _3121_ vssd1 vssd1 vccd1 vccd1 _3388_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ _3311_ _3314_ _3315_ _3318_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5520_ _1844_ _1848_ _1851_ _1854_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5451_ _1141_ _3490_ _1002_ _3493_ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4402_ _0738_ _0427_ _0740_ _0742_ _0744_ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__o2111a_1
X_5382_ _0563_ _0584_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__nand2_1
X_4333_ egd_top.BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7121_ _0071_ _0232_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7052_ _0002_ _0163_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_4264_ _0606_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6003_ _2332_ _2333_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ _3119_ _0484_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6905_ _3042_ _3043_ clknet_1_0__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6836_ _3024_ vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6767_ _2955_ _2960_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__or2_1
X_3979_ _0322_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__buf_2
X_5718_ _3497_ _0389_ _0701_ _0392_ _2050_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6698_ _2881_ _2894_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5649_ _1861_ _1982_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 la_data_in_47_32[15] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4951_ _1244_ _1260_ _1274_ _1289_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3902_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _3440_ sky130_fd_sc_hd__inv_2
X_4882_ _1209_ _1214_ _1218_ _1221_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6621_ _2817_ _2818_ vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__nand2_1
X_3833_ _3370_ vssd1 vssd1 vccd1 vccd1 _3371_ sky130_fd_sc_hd__buf_4
X_3764_ _3301_ _3214_ vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__nor2_4
XFILLER_0_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6552_ _2751_ _2752_ vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3695_ _3232_ egd_top.BitStream_buffer.pc\[2\] _3216_ vssd1 vssd1 vccd1 vccd1 _3233_
+ sky130_fd_sc_hd__and3_1
X_6483_ _3276_ _3090_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__nor2_1
X_5503_ _0437_ _0544_ _0743_ _0547_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5434_ _0679_ _3401_ _0840_ _3405_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7104_ _0054_ _0215_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
X_5365_ _3168_ _0464_ _3171_ _0468_ _1700_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__a221oi_1
X_5296_ _0569_ _3326_ _0564_ _3330_ _1631_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__a221oi_1
X_4316_ _0601_ _3332_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__o21ai_1
X_4247_ _0585_ _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__nand2_1
X_7035_ _3072_ _3073_ clknet_1_0__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__o21ai_2
X_4178_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__clkbuf_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6819_ _3009_ vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5150_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__o21ai_1
X_5081_ _1408_ _1410_ _1413_ _1418_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__and4_1
X_4101_ _0444_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__clkbuf_4
X_4032_ _0375_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__buf_2
X_5983_ _0488_ _0448_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4934_ _0679_ _3452_ _0840_ _3456_ _1272_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__a221oi_1
X_4865_ _1199_ _1201_ _1204_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__and3_1
XANTENNA_12 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6604_ _2783_ _2792_ vssd1 vssd1 vccd1 vccd1 _2802_ sky130_fd_sc_hd__nand2_1
XANTENNA_45 _3242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__clkbuf_4
X_4796_ _1134_ _1135_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__nand2_1
X_3747_ _3284_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__clkbuf_2
X_6535_ _2737_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3678_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__inv_2
X_6466_ _2693_ _2694_ _2695_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5417_ _1742_ _1746_ _1749_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__and4_1
X_6397_ net10 _0589_ _2619_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5348_ _0634_ _0390_ _0796_ _0393_ _1683_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__a221oi_1
X_5279_ _3237_ _3264_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__nand2_1
X_7018_ _3069_ _3070_ clknet_1_0__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_0__3077_ _3077_ vssd1 vssd1 vccd1 vccd1 clknet_0__3077_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4650_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3601_ _3092_ _3084_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__nand2_1
Xinput10 la_data_in_47_32[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_4
Xinput21 la_oenb_64 vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4581_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__inv_2
X_6320_ net3 _3340_ _2470_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__mux2_1
X_3532_ net37 net36 vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__nor2_1
X_6251_ _2546_ _2536_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__and2_1
X_5202_ _3508_ _3238_ _3511_ _3213_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6182_ _2499_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5133_ _0588_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _1471_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ _1400_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4015_ _3289_ _0344_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5966_ _0416_ _3195_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5897_ _3244_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _2228_
+ sky130_fd_sc_hd__nand2_1
X_4917_ _3386_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _1256_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4848_ _1174_ _1179_ _1183_ _1187_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__and4_1
X_4779_ _3386_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _1119_
+ sky130_fd_sc_hd__nand2_1
X_6518_ net13 _0916_ _2707_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6449_ _2682_ _2668_ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5820_ _0704_ _3489_ _3503_ _3492_ _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__o221a_1
X_5751_ _2079_ _2081_ _2083_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__and3_1
X_4702_ _0451_ _0435_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5682_ _0971_ _3423_ _2014_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _0971_ _3350_ _0973_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__o21ai_1
X_4564_ _0891_ _0897_ _0901_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6303_ _2582_ _2580_ vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6234_ net13 _0801_ _2516_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__mux2_1
X_4495_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6165_ _2487_ _3197_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__and2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _0503_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _1454_
+ sky130_fd_sc_hd__nand2_1
X_6096_ _0455_ _3152_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__nand2_1
X_5047_ _0823_ _3361_ _0972_ _3365_ _1384_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6998_ _3026_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__buf_4
X_5949_ _0337_ egd_top.BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _2280_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ _0623_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6921_ clknet_1_1__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__buf_1
X_6852_ _3025_ _3028_ clknet_1_0__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5803_ _3358_ _3400_ _3362_ _3404_ _2134_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__a221oi_1
X_6783_ _2844_ _2949_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__nor2_1
X_3995_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5734_ _2065_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5665_ _3334_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _1998_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4616_ _3270_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _0957_
+ sky130_fd_sc_hd__nand2_1
X_5596_ _1921_ _1924_ _1926_ _1929_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__and4_1
X_4547_ _0417_ _3152_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__nand2_1
X_4478_ _0786_ _3332_ _0819_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__o21ai_1
X_6217_ _2513_ _2523_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__and2_1
X_7197_ _0147_ _0308_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _2474_ _2475_ _2471_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__o21ai_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _0724_ _0366_ _2408_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3780_ _3317_ vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__buf_2
XFILLER_0_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5450_ _3496_ _0708_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4401_ _0743_ _0439_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__or2_1
X_5381_ _1712_ _1714_ _1716_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4332_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__buf_2
X_7120_ _0070_ _0231_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_7051_ _0001_ _0162_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[94\]
+ sky130_fd_sc_hd__dfxtp_1
X_4263_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6002_ _0587_ _0916_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4194_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6904_ _3042_ _3043_ clknet_1_0__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6835_ _3023_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__clkbuf_8
X_3978_ _3515_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__clkbuf_2
X_6766_ _2865_ _2956_ _2959_ vssd1 vssd1 vccd1 vccd1 _2960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5717_ _0693_ _0395_ _2049_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6697_ _2887_ _2893_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5648_ _3149_ _1981_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__nor2_1
X_5579_ _0327_ _3296_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__3074_ clknet_0__3074_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3074_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 la_data_in_47_32[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_4
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4950_ _1278_ _1280_ _1283_ _1288_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__and4_1
X_3901_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _3439_ sky130_fd_sc_hd__clkbuf_4
X_4881_ _0573_ _0614_ _0577_ _0618_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__a221oi_1
X_6620_ _2797_ _2784_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__nor2_2
X_3832_ _3369_ vssd1 vssd1 vccd1 vccd1 _3370_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6551_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1 vccd1
+ _2752_ sky130_fd_sc_hd__inv_2
X_3763_ _3276_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__nand2_8
X_5502_ _0452_ _0521_ _0746_ _0525_ _1836_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__a221oi_1
X_6482_ _2703_ _2693_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[2\] sky130_fd_sc_hd__xnor2_4
X_3694_ _3231_ vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5433_ _1644_ _3408_ _1767_ _3411_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__o22ai_1
X_5364_ _1698_ _1699_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__nand2_1
X_7103_ _0053_ _0214_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
X_4315_ _3335_ _0657_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__nand2_1
X_5295_ _1601_ _3332_ _1630_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4246_ _0588_ _0589_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__nand2_1
X_7034_ _3072_ _3073_ clknet_1_0__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__o21ai_2
X_4177_ _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__clkbuf_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6818_ _2993_ _2992_ _2814_ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__o21ai_1
X_6749_ _2872_ _2938_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5080_ _1414_ _1415_ _1416_ _1417_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__and4_1
X_4100_ _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4031_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5982_ _2295_ _2312_ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__nand2_1
X_4933_ _1270_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4864_ _0457_ _0537_ _0452_ _0541_ _1203_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6603_ _2775_ _2800_ vssd1 vssd1 vccd1 vccd1 _2801_ sky130_fd_sc_hd__nand2_2
XANTENNA_46 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3815_ _3352_ vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__buf_2
XANTENNA_24 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4795_ _3463_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _1135_
+ sky130_fd_sc_hd__nand2_1
X_3746_ _3283_ _3220_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__and2_1
X_6534_ _2736_ _3080_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6465_ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5416_ _0844_ _3305_ _0991_ _3310_ _1750_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3677_ _3214_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__inv_2
X_6396_ _2646_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
X_5347_ _0700_ _0396_ _1682_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5278_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__o21ai_1
X_7017_ _3069_ _3070_ clknet_1_0__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__o21ai_2
X_4229_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__buf_2
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _0768_ _0521_ _0919_ _0525_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__a221oi_1
Xinput11 la_data_in_47_32[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_4
Xinput22 la_oenb_65 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_1
X_3600_ net34 net33 vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__nand2_1
X_3531_ net35 vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6250_ net8 _3250_ _2515_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__mux2_1
X_5201_ _0649_ _3502_ _0810_ _3505_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6181_ _2498_ _2492_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__and2_4
X_5132_ _0583_ _1210_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__nand2_1
X_5063_ _3463_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1401_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4014_ _3174_ _0348_ _0352_ _0357_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5965_ _0411_ _3189_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5896_ _3236_ _0683_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__nand2_1
X_4916_ _0662_ _3361_ _0823_ _3365_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4847_ _0418_ _0464_ _0733_ _0468_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4778_ _3354_ _3361_ _0662_ _3365_ _1117_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a221oi_1
X_6517_ _2725_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
X_3729_ _3266_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__buf_4
X_6448_ net10 _0413_ net43 vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6379_ _2634_ _2624_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3059_ _3059_ vssd1 vssd1 vccd1 vccd1 clknet_0__3059_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5750_ _1039_ _0536_ _0461_ _0540_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4701_ _1037_ _0427_ _1038_ _1040_ _1041_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__o2111a_1
X_5681_ _3426_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _2014_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4632_ _3353_ _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4563_ _0413_ _0464_ _0731_ _0468_ _0904_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__a221oi_1
X_4494_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__buf_2
X_6302_ net8 _3428_ _2550_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__mux2_1
X_6233_ _2534_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ net4 _3497_ _2480_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__mux2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _0499_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _1453_
+ sky130_fd_sc_hd__nand2_1
X_6095_ _0450_ _3163_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5046_ _1382_ _3368_ _1383_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6997_ _3023_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__buf_4
X_5948_ _0332_ egd_top.BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _2279_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5879_ _0582_ _0916_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6920_ _3027_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6851_ _3025_ _3028_ clknet_1_0__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__o21ai_2
X_5802_ _3366_ _3407_ _0666_ _3410_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__o22ai_1
X_3994_ _0337_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__buf_4
X_6782_ _2973_ _2974_ _2818_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__nand3_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5733_ _0474_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _2066_
+ sky130_fd_sc_hd__nand2_1
X_5664_ _1987_ _1991_ _1994_ _1996_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4615_ _3263_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _0956_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5595_ _0947_ _0389_ _3497_ _0392_ _1928_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4546_ _0412_ _0418_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4477_ _3335_ _0818_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__nand2_1
X_6216_ net4 _3296_ _2516_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__mux2_1
X_7196_ _0146_ _0307_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ net45 _3124_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _0369_ _3208_ vssd1 vssd1 vccd1 vccd1 _2408_ sky130_fd_sc_hd__nand2_1
X_5029_ _0991_ _3254_ _1130_ _3258_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__inv_2
X_5380_ _0435_ _0537_ _0741_ _0541_ _1715_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4331_ _0660_ _0665_ _0669_ _0673_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7050_ _0000_ _0161_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_4262_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__buf_2
X_6001_ _0582_ _0518_ vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4193_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6903_ _3042_ _3043_ clknet_1_0__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6834_ net19 vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__buf_4
X_3977_ _3307_ _3469_ vssd1 vssd1 vccd1 vccd1 _3515_ sky130_fd_sc_hd__and2_1
X_6765_ _2958_ _2865_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5716_ _0398_ _0695_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__nand2_1
X_6696_ _2889_ _2892_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5647_ _1918_ _1979_ _1980_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__nand3_1
X_5578_ _0322_ _3238_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__nand2_1
X_4529_ _0857_ _0860_ _0864_ _0870_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__and4_1
X_7179_ _0129_ _0290_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 la_data_in_47_32[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_4
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3900_ _3437_ vssd1 vssd1 vccd1 vccd1 _3438_ sky130_fd_sc_hd__buf_2
X_4880_ _1082_ _0621_ _1219_ _0624_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__o22ai_1
X_3831_ _3283_ _3121_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3762_ egd_top.BitStream_buffer.BS_buffer\[26\] vssd1 vssd1 vccd1 vccd1 _3300_ sky130_fd_sc_hd__clkbuf_4
X_6550_ _2749_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__nand2_1
X_5501_ _1202_ _0528_ _1334_ _0531_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__o22ai_1
X_3693_ _3115_ _3230_ vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__nand2_2
X_6481_ _2694_ _2695_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__nand2_2
X_5432_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__inv_2
X_5363_ _0475_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _1699_
+ sky130_fd_sc_hd__nand2_1
X_7102_ _0052_ _0213_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_4314_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5294_ _3335_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _1630_
+ sky130_fd_sc_hd__nand2_1
X_4245_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__clkbuf_4
X_7033_ _3072_ _3073_ clknet_1_0__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__o21ai_2
X_4176_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6817_ _3005_ _2999_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6748_ _2872_ _2938_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6679_ _2872_ _2875_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3056_ clknet_0__3056_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3056_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4030_ _3251_ _0344_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5981_ _2299_ _2303_ _2307_ _2311_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__and4_1
X_4932_ _3463_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _1271_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6602_ _2797_ _2783_ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__nor2_1
X_4863_ _1065_ _0544_ _1202_ _0547_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__o22ai_1
XANTENNA_14 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _3351_ vssd1 vssd1 vccd1 vccd1 _3352_ sky130_fd_sc_hd__clkbuf_2
XANTENNA_36 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4794_ _3459_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _1134_
+ sky130_fd_sc_hd__nand2_1
X_6533_ net8 _0534_ _2706_ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__mux2_1
X_3745_ _3282_ vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__inv_2
X_6464_ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5415_ _1626_ _3314_ _3440_ _3318_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__o22ai_1
X_3676_ _3114_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6395_ _2644_ _2645_ vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__and2_1
X_5346_ _0399_ _0947_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__nand2_1
X_5277_ _1487_ _1613_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__nor2_1
X_7016_ _3069_ _3070_ clknet_1_0__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__o21ai_2
X_4228_ _0551_ _0556_ _0557_ _0560_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__a221oi_1
X_4159_ _0502_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput12 la_data_in_47_32[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_4
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput23 wb_rst_i vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_4
X_3530_ _3087_ _3088_ _3090_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a21oi_1
X_5200_ _0855_ _3490_ _0697_ _3493_ _1536_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__o221a_1
X_6180_ net14 _0339_ _2480_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5131_ _0589_ _0556_ _0584_ _0560_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__a221oi_1
X_5062_ _3459_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _1400_
+ sky130_fd_sc_hd__nand2_1
X_4013_ _0354_ egd_top.BitStream_buffer.BS_buffer\[118\] _0356_ egd_top.BitStream_buffer.BS_buffer\[119\]
+ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5964_ _2286_ _2289_ _2291_ _2294_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5895_ _3150_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__o21ai_1
X_4915_ _1252_ _3368_ _1253_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4846_ _1184_ _1185_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6516_ _2724_ _2689_ vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__and2_1
X_4777_ _1115_ _3368_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__o21ai_1
X_3728_ _3241_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__and3_1
X_6447_ _2681_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
X_3659_ _3200_ _3197_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__and2_1
X_6378_ net16 _0551_ _2620_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__mux2_1
X_5329_ _3508_ _3213_ _3511_ _3224_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4700_ _0738_ _0439_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__or2_1
X_5680_ _3372_ _3400_ _3358_ _3404_ _2012_ vssd1 vssd1 vccd1 vccd1 _2013_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4631_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__clkbuf_4
X_4562_ _0902_ _0903_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4493_ _0821_ _0826_ _0830_ _0834_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__and4_1
X_6301_ _2581_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_6232_ _2513_ _2533_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__and2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _2486_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__clkbuf_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _0920_ _0486_ _1451_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__o21ai_1
X_6094_ _0349_ _0426_ _2421_ _2422_ _2423_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__o2111a_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _3371_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _1383_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6996_ _3063_ _3064_ clknet_1_0__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__o21ai_2
X_5947_ _0327_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _2278_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5878_ _1073_ _0555_ _1210_ _0559_ _2209_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4829_ _3199_ _0390_ _3202_ _0393_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6850_ _3025_ _3028_ clknet_1_0__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6781_ _2943_ _2941_ _2971_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _2122_ _2125_ _2128_ _2132_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__and4_1
X_3993_ _0336_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5732_ _0470_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _2065_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ _1130_ _3304_ _3395_ _3309_ _1995_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4614_ _0801_ _3223_ _3300_ _3229_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5594_ _3468_ _0395_ _1927_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4545_ _0876_ _0880_ _0883_ _0886_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4476_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__buf_2
X_7195_ _0145_ _0306_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[119\]
+ sky130_fd_sc_hd__dfxtp_1
X_6215_ _2522_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ net44 net46 vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__nor2_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _0947_ _0347_ _2405_ _2406_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__a211oi_1
X_5028_ _1364_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6979_ _3060_ _3061_ clknet_1_1__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4330_ _3380_ _3379_ _3322_ _3383_ _0672_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__a221oi_1
X_4261_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6000_ _1210_ _0555_ _1055_ _0559_ _2330_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4192_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6902_ _3042_ _3043_ clknet_1_0__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6833_ _2869_ _3018_ _3016_ _2900_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__a22o_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3976_ _3506_ _3513_ vssd1 vssd1 vccd1 vccd1 _3514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6764_ _2924_ _2957_ vssd1 vssd1 vccd1 vccd1 _2958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5715_ _0329_ _0375_ _0334_ _0378_ _2047_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__a221oi_1
X_6695_ _2890_ _2891_ _2810_ vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__o21ai_1
X_5646_ _0632_ _0334_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__nand2_1
X_5577_ _1909_ _1910_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4528_ _0866_ _0867_ _0868_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__and4_1
X_4459_ egd_top.BitStream_buffer.BS_buffer\[25\] vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7178_ _0128_ _0289_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ sky130_fd_sc_hd__dfxtp_2
X_6129_ _0781_ _0595_ _0932_ _0599_ _2458_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__a221oi_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _3367_ vssd1 vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__buf_2
X_3761_ _3275_ _3281_ _3286_ _3287_ _3298_ vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5500_ _1828_ _1832_ _1833_ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__and4b_1
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6480_ _3216_ _3090_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__nor2_1
X_3692_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5431_ _1755_ _1758_ _1761_ _1765_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__and4_1
X_5362_ _0471_ _3163_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__nand2_1
X_4313_ _0643_ _0647_ _0652_ _0655_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__and4_1
X_7101_ _0051_ _0212_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_5293_ _1618_ _1622_ _1625_ _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__and4_1
X_7032_ _3072_ _3073_ clknet_1_0__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__o21ai_2
X_4244_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__buf_2
X_4175_ _3302_ _0484_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__and2_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6816_ _2927_ _3006_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__nor2_1
X_6747_ _2940_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _3497_ sky130_fd_sc_hd__clkbuf_4
X_6678_ _2873_ _2874_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__nand2_1
X_5629_ _0562_ _0577_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5980_ _3183_ _0463_ _3186_ _0467_ _2310_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4931_ _3459_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1270_
+ sky130_fd_sc_hd__nand2_1
X_4862_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6601_ _2797_ _2798_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__nor2_2
X_3813_ _3217_ _3121_ vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__and2_1
XANTENNA_26 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _0991_ _3435_ _3438_ _1130_ _1132_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_48 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3744_ _3277_ _3231_ vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6532_ _2735_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3675_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__clkbuf_4
X_6463_ _2691_ _3113_ _2692_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5414_ _0801_ _3281_ _3286_ _3300_ _1748_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6394_ net39 vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__buf_2
X_5345_ _3476_ _0376_ _3482_ _0379_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5276_ _3212_ _1612_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__nor2_1
X_7015_ _3069_ _3070_ clknet_1_0__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__o21ai_2
X_4227_ _0565_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__3074_ _3074_ vssd1 vssd1 vccd1 vccd1 clknet_0__3074_ sky130_fd_sc_hd__clkbuf_16
X_4158_ _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__clkbuf_2
X_4089_ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 la_data_in_47_32[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_4
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__3038_ clknet_0__3038_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3038_
+ sky130_fd_sc_hd__clkbuf_16
X_5130_ _1466_ _1467_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__nand2_1
X_5061_ _3395_ _3435_ _3438_ _3402_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__a221oi_1
X_4012_ _0355_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5963_ _0695_ _0389_ _3476_ _0392_ _2293_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4914_ _3371_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _1253_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5894_ _2105_ _2225_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4845_ _0475_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1185_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4776_ _3371_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _1116_
+ sky130_fd_sc_hd__nand2_1
X_3727_ _3263_ _3264_ vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6515_ net14 _0765_ _2707_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6446_ _2680_ _2668_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__and2_1
X_3658_ net10 _3199_ _3158_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__mux2_1
X_3589_ _3142_ _3144_ _3081_ _3145_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__o211a_1
X_6377_ _2633_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__clkbuf_1
X_5328_ _0810_ _3502_ _0960_ _3505_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__o22ai_1
X_5259_ _0584_ _0556_ _0573_ _0560_ _1595_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4630_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4561_ _0475_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _0903_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6300_ _2579_ _2580_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4492_ _3322_ _3379_ _3327_ _3383_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__a221oi_2
X_6231_ net14 _0639_ _2516_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _2485_ _3197_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__and2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _0489_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _1451_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _1022_ _0438_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__or2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6995_ _3063_ _3064_ clknet_1_1__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__o21ai_2
X_5946_ _0322_ _0639_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5877_ _2207_ _2208_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4828_ _0881_ _0396_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4759_ _0683_ _3254_ _0844_ _3258_ _1098_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a221oi_1
X_6429_ _2669_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3992_ _3312_ _3469_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__and2_1
X_6780_ _2970_ _2972_ vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5800_ _0551_ _3378_ _0557_ _3382_ _2131_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__a221oi_1
X_5731_ _0465_ _0444_ _0446_ _0413_ _2063_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5662_ _0684_ _3313_ _3406_ _3317_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__o22ai_1
X_4613_ _0952_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5593_ _0398_ _0701_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__nand2_1
X_4544_ _3192_ _0390_ _3195_ _0393_ _0885_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__a221oi_1
X_4475_ _0805_ _0809_ _0813_ _0816_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__and4_1
X_6214_ _2521_ _2513_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__and2_1
X_7194_ _0144_ _0305_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _3124_ _2471_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__or2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _0353_ _0701_ _0355_ _0695_ vssd1 vssd1 vccd1 vccd1 _2406_ sky130_fd_sc_hd__a22o_1
X_5027_ _3270_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _1365_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6978_ _3060_ _3061_ clknet_1_0__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5929_ _3444_ _0840_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4260_ _3283_ _0552_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__and2_1
X_4191_ _3251_ _0484_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__and2_1
X_6901_ _3042_ _3043_ clknet_1_0__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6832_ _3021_ _3022_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__nand2_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3975_ _3508_ _3509_ _3511_ _3512_ vssd1 vssd1 vccd1 vccd1 _3513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6763_ _2931_ _2862_ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__nor2_1
X_5714_ _3483_ _0381_ _0697_ _0384_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__o22ai_1
X_6694_ _2763_ _2841_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5645_ _1948_ _1978_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5576_ _3507_ egd_top.BitStream_buffer.BS_buffer\[24\] _3510_ _0801_ vssd1 vssd1
+ vccd1 vccd1 _1910_ sky130_fd_sc_hd__a22o_1
X_4527_ _0338_ _0334_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4458_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] _3081_ vssd1
+ vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__o21ai_1
X_7177_ _0127_ _0288_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_6128_ _1350_ _0602_ _2457_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__o21ai_1
X_4389_ _0412_ _0731_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__nand2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _3474_ _3246_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__3071_ clknet_0__3071_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3071_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3760_ _3288_ _3291_ _3297_ vssd1 vssd1 vccd1 vccd1 _3298_ sky130_fd_sc_hd__o21ai_1
X_3691_ _3228_ vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__buf_2
X_5430_ _0597_ _3379_ _0569_ _3383_ _1764_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _0894_ _0445_ _0447_ _1039_ _1696_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__a221oi_2
X_4312_ _3306_ _3305_ _3271_ _3310_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _0683_ _3305_ _0844_ _3310_ _1627_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__a221oi_1
X_7100_ _0050_ _0211_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
X_4243_ _0586_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__clkbuf_2
X_7031_ _3072_ _3073_ clknet_1_0__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__o21ai_2
X_4174_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6815_ _2863_ _2932_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6746_ _2756_ _2814_ _2939_ vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3958_ _3495_ vssd1 vssd1 vccd1 vccd1 _3496_ sky130_fd_sc_hd__buf_2
X_6677_ _2814_ _2748_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__nand2_1
X_3889_ _3426_ vssd1 vssd1 vccd1 vccd1 _3427_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5628_ _1957_ _1959_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5559_ _0822_ _3423_ _1892_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4930_ _1130_ _3435_ _3438_ _3395_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4861_ _0534_ _0521_ _0538_ _0525_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6600_ _2783_ _2775_ vssd1 vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__or2_1
X_3812_ _3349_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_27 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4792_ _0676_ _3442_ _1131_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__o21ai_1
XANTENNA_16 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _1205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3743_ _3280_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__clkbuf_4
X_6531_ _2734_ _3080_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__and2_1
XANTENNA_49 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3674_ _3149_ vssd1 vssd1 vccd1 vccd1 _3212_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6462_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5413_ _0814_ _3291_ _1747_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6393_ net11 _0615_ _2619_ vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5344_ _0858_ _0382_ _3468_ _0385_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__o22ai_1
X_5275_ _1547_ _1610_ _1611_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__nand3_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7014_ _3069_ _3070_ clknet_1_0__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__o21ai_2
X_4226_ _0568_ _0569_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4157_ _3289_ _0483_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__and2_1
X_4088_ _3217_ _0407_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6729_ _2902_ _2924_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 la_data_in_47_32[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_4
XFILLER_0_3_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ _0985_ _3442_ _1397_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__o21ai_1
X_4011_ _3226_ _0345_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5962_ _0697_ _0395_ _2292_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4913_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5893_ _3149_ _2224_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4844_ _0471_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _1184_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4775_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__inv_2
X_3726_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__clkbuf_4
X_6514_ _2723_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6445_ net11 _0465_ net43 vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__mux2_1
X_3657_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__buf_2
X_3588_ _3140_ _3141_ net33 vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__a21o_1
X_6376_ _2632_ _2624_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__and2_1
X_5327_ _1002_ _3490_ _0855_ _3493_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__o221a_1
X_5258_ _1593_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__3056_ _3056_ vssd1 vssd1 vccd1 vccd1 clknet_0__3056_ sky130_fd_sc_hd__clkbuf_16
X_5189_ _3402_ _3435_ _3438_ _0675_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__a221oi_1
X_4209_ _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4560_ _0471_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _0902_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4491_ _0831_ _0832_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6230_ _2532_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ net5 _0947_ _2480_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__mux2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _1432_ _1449_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _0433_ _3174_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__nand2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _3376_ _3343_ _3380_ _3347_ _1380_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6994_ _3063_ _3064_ clknet_1_1__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5945_ _2274_ _2275_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__nor2_1
X_5876_ _0567_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _2208_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4827_ _0399_ _3205_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4758_ _1096_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3709_ _3245_ _3246_ vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__nand2_1
X_4689_ _0724_ _0396_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__o21ai_1
X_6428_ _2667_ _2668_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6359_ net7 _0818_ _2620_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3991_ _0333_ _0334_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5730_ _2061_ _2062_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5661_ _3306_ _3280_ _3285_ _3271_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4612_ _3245_ _3224_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__nand2_1
X_5592_ _0339_ _0375_ _0329_ _0378_ _1925_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4543_ _0383_ _0396_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4474_ _3271_ _3305_ _3264_ _3310_ _0815_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__a221oi_1
X_6213_ net5 _0648_ _2516_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__mux2_1
X_7193_ _0143_ _0304_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _2470_ _2472_ _3090_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a21oi_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6075_ _0700_ _0350_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__nor2_1
X_5026_ _3263_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _1364_
+ sky130_fd_sc_hd__nand2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6977_ _3060_ _3061_ clknet_1_1__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__o21ai_2
X_5928_ _0972_ _3416_ _3376_ _3420_ _2258_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5859_ _2178_ _2182_ _2186_ _2190_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4190_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6900_ _3042_ _3043_ clknet_1_0__leaf__3044_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__o21ai_2
X_6831_ _2999_ _2900_ vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__nand2_1
X_6762_ _2896_ _2927_ vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__nand2_1
X_3974_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _3512_ sky130_fd_sc_hd__buf_2
X_6693_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _2842_ vssd1 vssd1
+ vccd1 vccd1 _2890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5713_ _3202_ _0360_ _3205_ _0363_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5644_ _1962_ _1977_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5575_ _1100_ _3501_ _1237_ _3504_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4526_ _0333_ _0708_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__nand2_1
X_4457_ _0638_ _0799_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7176_ _0126_ _0287_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_6127_ _0605_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _2457_
+ sky130_fd_sc_hd__nand2_1
X_4388_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__clkbuf_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _2377_ _2380_ _2383_ _2387_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__and4_1
X_5009_ _1346_ _0603_ _1347_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3690_ _3227_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5360_ _1694_ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__nand2_1
X_4311_ _3315_ _3314_ _0653_ _3318_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__o22ai_1
X_5291_ _1499_ _3314_ _1626_ _3318_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4242_ _3267_ _0552_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__and2_1
X_7030_ _3072_ _3073_ clknet_1_1__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__o21ai_2
X_4173_ _0491_ _0506_ _0511_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__and4b_1
XFILLER_0_77_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6814_ _2986_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6745_ _2814_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1
+ vccd1 _2939_ sky130_fd_sc_hd__nand2_1
X_3957_ _3494_ vssd1 vssd1 vccd1 vccd1 _3495_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6676_ _2833_ _2752_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__nand2_1
X_3888_ _3425_ vssd1 vssd1 vccd1 vccd1 _3426_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5627_ _0894_ _0536_ _1039_ _0540_ _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5558_ _3426_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _1892_
+ sky130_fd_sc_hd__nand2_1
X_4509_ _3414_ _3452_ _3418_ _3456_ _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__a221oi_1
X_5489_ _3171_ _0464_ _3174_ _0468_ _1823_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__a221oi_1
X_7159_ _0109_ _0270_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3053_ clknet_0__3053_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3053_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4860_ _0542_ _0528_ _0545_ _0531_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__o22ai_1
X_3811_ _3226_ _3323_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__nand2_2
X_4791_ _3445_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _1131_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6530_ net9 _0919_ _2706_ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__mux2_1
XANTENNA_28 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _3242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3742_ _3279_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3673_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] _3081_ vssd1
+ vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__o21ai_1
X_6461_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__nor2_1
X_5412_ _3295_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _1747_
+ sky130_fd_sc_hd__nand2_1
X_6392_ _2643_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5343_ _3192_ _0361_ _3195_ _0364_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5274_ _0633_ _3482_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nand2_1
X_7013_ _3069_ _3070_ clknet_1_1__leaf__3071_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__o21ai_2
X_4225_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__clkbuf_4
X_4156_ _0499_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _0500_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4087_ _0430_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _0431_
+ sky130_fd_sc_hd__nand2_1
X_4989_ _1192_ _0494_ _0496_ _0510_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__a221oi_1
X_6728_ _2913_ _2923_ _2740_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6659_ _2799_ _2856_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput15 la_data_in_47_32[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4010_ _0353_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__buf_2
X_5961_ _0398_ _3482_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4912_ _0972_ _3343_ _3376_ _3347_ _1250_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_87_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5892_ _2162_ _2222_ _2223_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__nand3_1
X_4843_ _0746_ _0445_ _0447_ _0739_ _1182_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _0823_ _3343_ _0972_ _3347_ _1113_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3725_ _3262_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__buf_2
X_6513_ _2722_ _2689_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6444_ _2679_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3656_ _3198_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3587_ _3102_ _3104_ vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__nor2_1
X_6375_ net2 _0564_ _2620_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__mux2_1
X_5326_ _3496_ _0324_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5257_ _0568_ _0615_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__nand2_1
X_4208_ _3396_ _3218_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _0552_
+ sky130_fd_sc_hd__and3_2
X_5188_ _1124_ _3442_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__o21ai_1
X_4139_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4490_ _3390_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _0832_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ _2484_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _1436_ _1440_ _1444_ _1448_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__and4_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _0429_ _3168_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__nand2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _1378_ _3350_ _1379_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6993_ _3063_ _3064_ clknet_1_1__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__o21ai_2
X_5944_ _3507_ egd_top.BitStream_buffer.BS_buffer\[27\] _3510_ egd_top.BitStream_buffer.BS_buffer\[28\]
+ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5875_ _0562_ _0932_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4826_ _0947_ _0376_ _3497_ _0379_ _1165_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4757_ _3270_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _1097_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3708_ egd_top.BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4688_ _0399_ _3202_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nand2_1
X_6427_ _3079_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__clkbuf_2
X_3639_ _3185_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6358_ _2619_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__clkbuf_4
X_5309_ _1518_ _3408_ _1644_ _3411_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__o22ai_1
X_6289_ net12 _3449_ _2550_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3038_ _3038_ vssd1 vssd1 vccd1 vccd1 clknet_0__3038_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 net48 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5660_ _1104_ _3290_ _1992_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__o21ai_1
X_4611_ _3237_ _0639_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5591_ _0693_ _0381_ _3483_ _0384_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__o22ai_1
X_4542_ _0399_ _3199_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__nand2_1
X_4473_ _0653_ _3314_ _0814_ _3318_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6212_ _2520_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
X_7192_ _0142_ _0303_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _2471_ egd_top.BitStream_buffer.buffer_index\[5\] egd_top.BitStream_buffer.buffer_index\[4\]
+ _3132_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__a31o_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6074_ _2361_ _2375_ _2388_ _2403_ vssd1 vssd1 vccd1 vccd1 _2404_ sky130_fd_sc_hd__and4_1
X_5025_ _3271_ _3223_ _3264_ _3229_ _1362_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__a221oi_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6976_ _3060_ _3061_ clknet_1_1__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__o21ai_2
X_5927_ _1248_ _3423_ _2257_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5858_ _3180_ _0463_ _3183_ _0467_ _2189_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__a221oi_1
X_4809_ _1147_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__nor2_1
X_5789_ _0941_ _3122_ _2120_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6830_ _3020_ _2869_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__nand2_1
X_6761_ _2954_ vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _3510_ vssd1 vssd1 vccd1 vccd1 _3511_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5712_ _0394_ _0366_ _2044_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__o21ai_1
X_6692_ _2788_ _2888_ _2799_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5643_ _1966_ _1970_ _1973_ _1976_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__and4_1
X_5574_ _3500_ _3489_ _1141_ _3492_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4525_ _0328_ _0324_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4456_ _3212_ _0798_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nor2_1
X_7175_ _0125_ _0286_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_4387_ _0719_ _0723_ _0726_ _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__and4_1
X_6126_ _0768_ _0575_ _0919_ _0579_ _2455_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__a221oi_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _0823_ _3451_ _0972_ _3455_ _2386_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__a221oi_1
X_5008_ _0606_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _1347_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6959_ _3026_ vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__buf_4
XFILLER_0_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5290_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__inv_2
X_4310_ egd_top.BitStream_buffer.BS_buffer\[26\] vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _0583_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__nand2_1
X_4172_ _0514_ _0515_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6813_ _3003_ _3004_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__nand2_1
X_6744_ _2875_ _2911_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3956_ _3292_ _3470_ vssd1 vssd1 vccd1 vccd1 _3494_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6675_ _2817_ _2831_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__nand2_2
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5626_ _0743_ _0543_ _0425_ _0546_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3887_ _3251_ _3397_ vssd1 vssd1 vccd1 vccd1 _3425_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5557_ _0840_ _3400_ _3372_ _3404_ _1890_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__a221oi_1
X_4508_ _0848_ _0849_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__nand2_1
X_5488_ _1821_ _1822_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4439_ _0583_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _0782_
+ sky130_fd_sc_hd__nand2_1
X_7158_ _0108_ _0269_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_6109_ _2437_ _2438_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__nand2_1
X_7089_ _0039_ _0200_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4790_ egd_top.BitStream_buffer.BS_buffer\[37\] vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__clkbuf_4
X_3810_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__inv_2
X_3741_ _3278_ _3220_ vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__and2_1
XANTENNA_29 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ _2690_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
X_3672_ _3210_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
X_5411_ _3402_ _3254_ _0675_ _3258_ _1745_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__a221oi_1
X_6391_ _2642_ _2624_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__and2_1
X_5342_ _1018_ _0367_ _1677_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5273_ _1577_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__nor2_1
X_7012_ clknet_1_0__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3071_ sky130_fd_sc_hd__buf_1
Xclkbuf_0__3071_ _3071_ vssd1 vssd1 vccd1 vccd1 clknet_0__3071_ sky130_fd_sc_hd__clkbuf_16
X_4224_ _0567_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__buf_2
X_4155_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4086_ _0429_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4988_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6727_ _2916_ _2919_ _2922_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__and3_1
X_3939_ _3475_ _3476_ vssd1 vssd1 vccd1 vccd1 _3477_ sky130_fd_sc_hd__nand2_1
X_6658_ _2787_ _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5609_ _0470_ _3171_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2_1
X_6589_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] _2787_ vssd1 vssd1 vccd1
+ vccd1 _2788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 la_data_in_47_32[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__3035_ clknet_0__3035_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3035_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5960_ _0324_ _0375_ _0708_ _0378_ _2290_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__a221oi_1
X_4911_ _1248_ _3350_ _1249_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__o21ai_1
X_5891_ _0632_ _0708_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _1180_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _1111_ _3350_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__o21ai_1
X_3724_ _3261_ vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__clkbuf_2
X_6512_ net15 _0515_ _2707_ vssd1 vssd1 vccd1 vccd1 _2722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6443_ _2678_ _2668_ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__and2_1
X_3655_ _3196_ _3197_ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3586_ _3105_ _3142_ _3081_ _3143_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6374_ _2631_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5325_ _3503_ _3472_ _1658_ _1659_ _1660_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__o2111a_1
X_5256_ _0563_ _0589_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__clkbuf_4
X_5187_ _3445_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _1524_
+ sky130_fd_sc_hd__nand2_1
X_4138_ egd_top.BitStream_buffer.pc\[5\] _3120_ _3396_ vssd1 vssd1 vccd1 vccd1 _0482_
+ sky130_fd_sc_hd__or3_2
X_4069_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _3152_ _0464_ _3163_ _0468_ _1447_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__a221oi_1
X_6090_ _0383_ _0408_ _2417_ _2418_ _2419_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _3353_ _3322_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__nand2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6992_ _3063_ _3064_ clknet_1_0__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5943_ _3315_ _3501_ _0653_ _3504_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__o22ai_1
X_5874_ _2201_ _2203_ _2205_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4825_ _1026_ _0382_ _3491_ _0385_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _3263_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _1096_
+ sky130_fd_sc_hd__nand2_1
X_3707_ _3244_ vssd1 vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__buf_2
X_4687_ _0796_ _0376_ _0947_ _0379_ _1027_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_3_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6426_ net2 _0739_ _2656_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__mux2_1
X_3638_ _3184_ _3166_ vssd1 vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6357_ _2471_ _3126_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__nand2_4
X_3569_ egd_top.BitStream_buffer.pc\[6\] _3108_ _3123_ _3126_ vssd1 vssd1 vccd1 vccd1
+ _3127_ sky130_fd_sc_hd__or4b_1
X_5308_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__inv_2
X_6288_ _2572_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
X_5239_ _1563_ _1567_ _1571_ _1575_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 _2655_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_2
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4610_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] _3081_ vssd1
+ vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__o21ai_1
X_5590_ _3199_ _0360_ _3202_ _0363_ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4541_ _0634_ _0376_ _0796_ _0379_ _0882_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4472_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6211_ _2519_ _2513_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__and2_1
X_7191_ _0141_ _0302_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[123\]
+ sky130_fd_sc_hd__dfxtp_1
X_6142_ _3156_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__buf_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__3077_ clknet_0__3077_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3077_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _2392_ _2394_ _2397_ _2402_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__and4_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _1360_ _1361_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__nand2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6975_ _3060_ _3061_ clknet_1_1__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__o21ai_2
X_5926_ _3426_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _2257_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5857_ _2187_ _2188_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__nand2_1
X_4808_ _3508_ _0648_ _3511_ _3296_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a22o_1
X_5788_ _3334_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _2120_
+ sky130_fd_sc_hd__nand2_1
X_4739_ _1078_ _0603_ _1079_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6409_ _2471_ net42 _2475_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__nand3_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6760_ _2945_ _2953_ _2740_ vssd1 vssd1 vccd1 vccd1 _2954_ sky130_fd_sc_hd__a21oi_2
X_3972_ _3119_ _3470_ vssd1 vssd1 vccd1 vccd1 _3510_ sky130_fd_sc_hd__and2_2
X_5711_ _0369_ _3199_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__nand2_1
X_6691_ _2756_ _2786_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__nor2_1
X_5642_ _1055_ _0613_ _1192_ _0617_ _1975_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5573_ _3495_ _0865_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4524_ _0323_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4455_ _0715_ _0795_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__nand3_2
X_7174_ _0124_ _0285_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4386_ _3189_ _0390_ _3192_ _0393_ _0728_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a221oi_1
X_6125_ _2453_ _2454_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__nand2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _2384_ _2385_ vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__nand2_1
X_5007_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6958_ _3023_ vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__buf_4
X_5909_ _2230_ _2234_ _2237_ _2239_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__and4_1
X_6889_ _3039_ _3040_ clknet_1_1__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4240_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__clkbuf_4
X_4171_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6812_ _2981_ _2900_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3955_ _3492_ vssd1 vssd1 vccd1 vccd1 _3493_ sky130_fd_sc_hd__buf_2
X_6743_ _2930_ _2933_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__nand2_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6674_ _2826_ _2870_ _2871_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__nand3b_2
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5625_ _0746_ _0520_ _0739_ _0524_ _1958_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__a221oi_1
X_3886_ _3423_ vssd1 vssd1 vccd1 vccd1 _3424_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5556_ _1767_ _3407_ _3422_ _3410_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__o22ai_1
X_4507_ _3463_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _0849_
+ sky130_fd_sc_hd__nand2_1
X_5487_ _0475_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _1822_
+ sky130_fd_sc_hd__nand2_1
X_4438_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7157_ _0107_ _0268_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_4369_ _0338_ _0329_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__nand2_1
X_6108_ _0502_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _2438_
+ sky130_fd_sc_hd__nand2_1
X_7088_ _0038_ _0199_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _1506_ _3367_ _2368_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3740_ _3277_ _3240_ vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__nor2_8
XANTENNA_19 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3671_ _3209_ _3197_ vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__and2_1
X_5410_ _1743_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__nand2_1
X_6390_ net12 _0611_ _2619_ vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5341_ _0370_ _3189_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7011_ _3026_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__buf_4
X_5272_ _1592_ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__nand2_1
X_4223_ _0566_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__clkbuf_2
X_4154_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__clkbuf_2
X_4085_ _0428_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6726_ _2920_ _2921_ _2801_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__a21o_1
X_4987_ _0503_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _1326_
+ sky130_fd_sc_hd__nand2_1
X_3938_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _3476_ sky130_fd_sc_hd__clkbuf_4
X_6657_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3869_ _3242_ _3398_ vssd1 vssd1 vccd1 vccd1 _3407_ sky130_fd_sc_hd__nand2_2
X_6588_ _2786_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5608_ _0461_ _0444_ _0446_ _0465_ _1941_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__a221oi_1
X_5539_ _3440_ _3313_ _0684_ _3317_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__o22ai_1
X_7209_ _0159_ _0320_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput17 la_data_in_49_48[0] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4910_ _3353_ _3380_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__nand2_1
X_5890_ _2192_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _0456_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _1181_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4772_ _3353_ _3376_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3723_ _3260_ _3219_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__and2_1
X_6511_ _2721_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6442_ net12 _0461_ net43 vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__mux2_1
X_3654_ _3165_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__buf_8
XFILLER_0_70_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3585_ _3142_ _3101_ vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__nand2_1
X_6373_ _2630_ _2624_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__and2_1
X_5324_ _0861_ _3485_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5255_ _1586_ _1588_ _1591_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__and3_1
Xclkbuf_0__3053_ _3053_ vssd1 vssd1 vccd1 vccd1 clknet_0__3053_ sky130_fd_sc_hd__clkbuf_16
X_4206_ _0517_ _0533_ _0549_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5186_ _3362_ _3417_ _3340_ _3421_ _1522_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__a221oi_1
X_4137_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ _0411_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6709_ _2814_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1
+ vccd1 _2905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5040_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6991_ _3063_ _3064_ clknet_1_1__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__o21ai_2
X_5942_ _0861_ _3489_ _0704_ _3492_ _2272_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5873_ _0461_ _0536_ _0465_ _0540_ _2204_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4824_ _3180_ _0361_ _3183_ _0364_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4755_ _3300_ _3223_ _3306_ _3229_ _1094_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _3243_ vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4686_ _0881_ _0382_ _1026_ _0385_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__o22ai_1
X_6425_ _2666_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3637_ net15 _3183_ _3159_ vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3568_ _3124_ _3125_ net47 vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__and3_1
X_6356_ _2618_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5307_ _1632_ _1635_ _1638_ _1642_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__and4_1
X_6287_ _2571_ _2559_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__and2_1
X_5238_ _3163_ _0464_ _3168_ _0468_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__a221oi_1
X_5169_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 egd_top.BitStream_buffer.buffer_index\[5\] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4540_ _0724_ _0382_ _0881_ _0385_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__o22ai_1
X_4471_ _0648_ _3281_ _3286_ _3296_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6210_ net6 _3287_ _2516_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7190_ _0140_ _0301_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[124\]
+ sky130_fd_sc_hd__dfxtp_1
X_6141_ _2469_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__clkbuf_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _2398_ _2399_ _2400_ _2401_ vssd1 vssd1 vccd1 vccd1 _2402_ sky130_fd_sc_hd__and4_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _3245_ _3300_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__nand2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6974_ _3060_ _3061_ clknet_1_1__leaf__3062_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _3362_ _3400_ _3340_ _3404_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5856_ _0474_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _2188_
+ sky130_fd_sc_hd__nand2_1
X_4807_ _1007_ _3502_ _1146_ _3505_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5787_ _2109_ _2113_ _2116_ _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__and4_1
X_4738_ _0606_ _0569_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4669_ _1008_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6408_ _2654_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_6339_ net12 _3376_ _2469_ vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3971_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _3509_ sky130_fd_sc_hd__clkbuf_4
X_5710_ _3208_ _0347_ _2041_ _2042_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__a211oi_1
X_6690_ _2884_ _2886_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__nand2_1
X_5641_ _1852_ _0620_ _1974_ _0623_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5572_ _0861_ _3471_ _1903_ _1904_ _1905_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__o2111a_1
X_4523_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4454_ _0633_ _0796_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7173_ _0123_ _0284_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4385_ _0380_ _0396_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_0__f__3059_ clknet_0__3059_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3059_
+ sky130_fd_sc_hd__clkbuf_16
X_6124_ _0587_ _0518_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__nand2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _3462_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _2385_
+ sky130_fd_sc_hd__nand2_1
X_5006_ _1210_ _0576_ _1055_ _0580_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__a221oi_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _3054_ _3055_ clknet_1_1__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__o21ai_2
X_5908_ _3402_ _3304_ _0675_ _3309_ _2238_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__a221oi_1
X_6888_ _3039_ _3040_ clknet_1_0__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5839_ _0398_ _3476_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__buf_2
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6811_ _3001_ _3002_ _2869_ vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__nand3_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3954_ _3283_ _3470_ vssd1 vssd1 vccd1 vccd1 _3492_ sky130_fd_sc_hd__nand2_2
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6742_ _2935_ _2937_ vssd1 vssd1 vccd1 vccd1 egd_top.exp_golomb_decoding.te_range\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6673_ net18 _3110_ _2864_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__or3_1
X_3885_ _3119_ _3398_ vssd1 vssd1 vccd1 vccd1 _3423_ sky130_fd_sc_hd__nand2_2
X_5624_ _1334_ _0527_ _1462_ _0530_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__o22ai_1
X_5555_ _1878_ _1881_ _1884_ _1888_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4506_ _3459_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _0848_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5486_ _0471_ _3168_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__nand2_1
X_4437_ _0557_ _0556_ _0776_ _0560_ _0779_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__a221oi_1
X_7156_ _0106_ _0267_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6107_ _0498_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _2437_
+ sky130_fd_sc_hd__nand2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _0333_ _0324_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__nand2_1
X_4299_ _0640_ _0641_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__nand2_1
X_7087_ _0037_ _0198_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ _3370_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _2368_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3050_ clknet_0__3050_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3050_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3670_ net1 _3208_ _3158_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5340_ _3199_ _0348_ _1674_ _1675_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__a211oi_1
X_5271_ _1596_ _1600_ _1604_ _1607_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__and4_1
X_4222_ _3242_ _0552_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__and2_1
X_7010_ _3023_ vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__clkbuf_8
X_4153_ _3292_ _0483_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ _3242_ _0406_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4986_ _0499_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _1325_
+ sky130_fd_sc_hd__nand2_1
X_3937_ _3474_ vssd1 vssd1 vccd1 vccd1 _3475_ sky130_fd_sc_hd__buf_2
X_6725_ _2882_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] vssd1 vssd1
+ vccd1 vccd1 _2921_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3868_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _3406_ sky130_fd_sc_hd__inv_2
X_6656_ _2853_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__inv_2
X_6587_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__nor2_1
X_5607_ _1939_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__nand2_1
X_3799_ _3335_ _3336_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__nand2_1
X_5538_ _3300_ _3280_ _3285_ _3306_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__a221oi_1
X_7208_ _0158_ _0319_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dfxtp_2
X_5469_ _3482_ _0376_ _0339_ _0379_ _1803_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__a221oi_1
X_7139_ _0089_ _0250_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 la_data_in_49_48[1] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4840_ _0451_ _0741_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__nand2_1
X_6510_ _2720_ _2689_ vssd1 vssd1 vccd1 vccd1 _2721_ sky130_fd_sc_hd__and2_1
X_4771_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__inv_2
X_3722_ _3259_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6441_ _2677_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
X_3653_ net11 _3195_ _3158_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__mux2_1
X_6372_ net3 _0569_ _2620_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__mux2_1
X_3584_ _3140_ _3141_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__nand2_1
X_5323_ _3480_ _0708_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5254_ _0739_ _0537_ _0435_ _0541_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__a221oi_1
X_4205_ _0534_ _0537_ _0538_ _0541_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__a221oi_1
X_5185_ _1382_ _3424_ _1521_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _0403_ _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nand2_1
X_4067_ _0410_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6708_ _2833_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1
+ vccd1 _2904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6639_ _2836_ _2817_ vssd1 vssd1 vccd1 vccd1 _2837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6990_ _3063_ _3064_ clknet_1_1__leaf__3065_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__o21ai_2
X_5941_ _3495_ _3275_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5872_ _0738_ _0543_ _0892_ _0546_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4823_ _1161_ _0367_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4754_ _1092_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__nand2_1
X_3705_ _3242_ _3219_ vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4685_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__inv_2
X_6424_ _2665_ _2645_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__and2_1
X_3636_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3567_ egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 _3125_
+ sky130_fd_sc_hd__inv_2
X_6355_ _2617_ _2601_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__and2_1
X_6286_ net13 _0836_ _2551_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5306_ _0593_ _3379_ _0597_ _3383_ _1641_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5237_ _1572_ _1573_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__3035_ _3035_ vssd1 vssd1 vccd1 vccd1 clknet_0__3035_ sky130_fd_sc_hd__clkbuf_16
X_5168_ _0597_ _3326_ _0569_ _3330_ _1504_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__a221oi_1
X_5099_ _0430_ _0461_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__nand2_1
X_4119_ _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold7 egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4470_ _0810_ _3291_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6140_ _2468_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__buf_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _0337_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _2401_
+ sky130_fd_sc_hd__nand2_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _3237_ _3306_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__nand2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6973_ clknet_1_1__leaf__3030_ vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__buf_1
XFILLER_0_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _0666_ _3407_ _0827_ _3410_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5855_ _0470_ _3177_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4806_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5786_ _3395_ _3304_ _3402_ _3309_ _2117_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4737_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__inv_2
X_4668_ _3508_ _3287_ _3511_ _0648_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6407_ _2653_ _2645_ vssd1 vssd1 vccd1 vccd1 _2654_ sky130_fd_sc_hd__and2_1
X_3619_ _3170_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__clkbuf_1
X_4599_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__inv_2
X_6338_ _2606_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__clkbuf_1
X_6269_ _2558_ _2559_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _3507_ vssd1 vssd1 vccd1 vccd1 _3508_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5640_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5571_ _1146_ _3484_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4522_ _0862_ _0863_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__nor2_1
X_4453_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7172_ _0122_ _0283_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4384_ _0399_ _3195_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__nand2_1
X_6123_ _0582_ _0522_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__nand2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _3458_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _2384_
+ sky130_fd_sc_hd__nand2_1
X_5005_ _1342_ _1343_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__nand2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6956_ _3054_ _3055_ clknet_1_1__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5907_ _3409_ _3313_ _0676_ _3317_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__o22ai_1
X_6887_ _3039_ _3040_ clknet_1_1__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__o21ai_2
X_5838_ _0334_ _0375_ _0324_ _0378_ _2169_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5769_ _0632_ _0324_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6810_ _2987_ _2988_ _2999_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__nand3_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6741_ _2936_ _2742_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3953_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _3491_ sky130_fd_sc_hd__inv_2
X_6672_ _2863_ _2868_ _2869_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3884_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _3422_ sky130_fd_sc_hd__inv_2
X_5623_ _1950_ _1954_ _1955_ _1956_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__and4b_1
XFILLER_0_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5554_ _0569_ _3378_ _0564_ _3382_ _1887_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4505_ _0683_ _3435_ _3438_ _0844_ _0846_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5485_ _1039_ _0445_ _0447_ _0461_ _1819_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4436_ _0777_ _0778_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__nand2_1
X_7155_ _0105_ _0266_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_4367_ _0328_ _0334_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6106_ _1462_ _0485_ _2435_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__o21ai_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _3245_ _3238_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__nand2_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _0036_ _0197_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ _0593_ _3342_ _0597_ _3346_ _2366_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6939_ _3051_ _3052_ clknet_1_0__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__o21ai_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5270_ _0932_ _0614_ _1073_ _0618_ _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4221_ _0563_ _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nand2_1
X_4152_ _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__buf_2
X_4083_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4985_ _0769_ _0486_ _1323_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3936_ _3473_ vssd1 vssd1 vccd1 vccd1 _3474_ sky130_fd_sc_hd__clkbuf_2
X_6724_ _2847_ _2841_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6655_ _2801_ _2850_ _2852_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__o21ai_1
X_3867_ _3404_ vssd1 vssd1 vccd1 vccd1 _3405_ sky130_fd_sc_hd__buf_2
X_6586_ _2785_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ sky130_fd_sc_hd__inv_2
X_5606_ _0455_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1940_
+ sky130_fd_sc_hd__nand2_1
X_3798_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__clkbuf_4
X_5537_ _0964_ _3290_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7207_ _0157_ _0318_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__dfxtp_2
X_5468_ _3468_ _0382_ _0693_ _0385_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__o22ai_1
X_4419_ _0760_ _0761_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__nand2_1
X_5399_ _0633_ _0339_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__nand2_1
X_7138_ _0088_ _0249_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_7069_ _0019_ _0180_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__3032_ clknet_0__3032_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3032_
+ sky130_fd_sc_hd__clkbuf_16
Xinput19 la_data_in_64 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _0818_ _3326_ _0607_ _3330_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_70_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3721_ _3232_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__and3_1
X_6440_ _2676_ _2668_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__and2_1
X_3652_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__clkbuf_4
X_3583_ _3082_ _3091_ net38 net36 vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__and4_1
X_6371_ _2629_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5322_ _3475_ _3509_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__nand2_1
X_5253_ _1462_ _0544_ _1589_ _0547_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__o22ai_1
X_4204_ _0542_ _0544_ _0545_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__o22ai_1
X_5184_ _3427_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _1521_
+ sky130_fd_sc_hd__nand2_1
X_4135_ _0424_ _0441_ _0460_ _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4066_ _3267_ _0407_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4968_ _1161_ _0409_ _1304_ _1305_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4899_ _3295_ _0639_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2_1
X_6707_ _2872_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__inv_2
X_3919_ _3316_ _3397_ vssd1 vssd1 vccd1 vccd1 _3457_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6638_ _2834_ _2835_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__nand2_1
X_6569_ _2762_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5940_ _3288_ _3471_ _2268_ _2269_ _2270_ vssd1 vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5871_ _0435_ _0520_ _0741_ _0524_ _2202_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4822_ _0370_ _3177_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__nand2_1
X_4753_ _3245_ _0639_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3704_ _3241_ egd_top.BitStream_buffer.pc\[2\] _3216_ vssd1 vssd1 vccd1 vccd1 _3242_
+ sky130_fd_sc_hd__and3_4
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6423_ net3 _0746_ _2656_ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4684_ _3177_ _0361_ _3180_ _0364_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__a221oi_1
X_3635_ _3182_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__clkbuf_1
X_3566_ net44 vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__inv_2
X_6354_ net1 _0657_ _2469_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__mux2_1
X_6285_ _2570_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
X_5305_ _1639_ _1640_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__nand2_1
X_5236_ _0475_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1573_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5167_ _1474_ _3332_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4118_ _3302_ _0407_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__and2_1
X_5098_ _0349_ _0409_ _1433_ _1434_ _1435_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4049_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold8 _3125_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__3074_ clknet_0__3074_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3074_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _0332_ egd_top.BitStream_buffer.BS_buffer\[24\] vssd1 vssd1 vccd1 vccd1 _2400_
+ sky130_fd_sc_hd__nand2_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__o21ai_1
X_6972_ _3026_ vssd1 vssd1 vccd1 vccd1 _3061_ sky130_fd_sc_hd__buf_4
X_5923_ _2243_ _2246_ _2249_ _2253_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5854_ _0413_ _0444_ _0446_ _0731_ _2185_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4805_ _0693_ _3490_ _3468_ _3493_ _1144_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5785_ _3406_ _3313_ _3409_ _3317_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__o22ai_1
X_4736_ _0932_ _0576_ _1073_ _0580_ _1076_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4667_ _0861_ _3502_ _1007_ _3505_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6406_ net1 _0577_ _2619_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__mux2_1
X_3618_ _3169_ _3166_ vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__and2_1
X_4598_ _0569_ _0596_ _0564_ _0600_ _0939_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__a221oi_1
X_6337_ _2605_ _2601_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__and2_1
X_3549_ net34 _3106_ vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__nor2_1
X_6268_ net39 vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__clkbuf_2
X_6199_ _2492_ _2510_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__and2_1
X_5219_ _0399_ _0796_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5570_ _3479_ _3509_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4521_ _3508_ _3275_ _3511_ _3287_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4452_ _0756_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__nor2_1
X_7171_ _0121_ _0282_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4383_ _3208_ _0376_ _0634_ _0379_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__a221oi_1
X_6122_ _1055_ _0555_ _1192_ _0559_ _2451_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__a221oi_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _3428_ _3434_ _3437_ _0679_ _2382_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__a221oi_1
X_5004_ _0588_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _1343_
+ sky130_fd_sc_hd__nand2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6955_ _3054_ _3055_ clknet_1_1__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__o21ai_2
X_5906_ _3264_ _3280_ _3285_ _3250_ _2236_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6886_ _3039_ _3040_ clknet_1_0__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5837_ _0697_ _0381_ _0855_ _0384_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5768_ _2070_ _2100_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__nor2_1
X_4719_ _0509_ _0916_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__nand2_1
X_5699_ _3507_ egd_top.BitStream_buffer.BS_buffer\[25\] _3510_ _3300_ vssd1 vssd1
+ vccd1 vccd1 _2032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ _2930_ _2934_ _2933_ vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__nand3_1
X_3952_ _3489_ vssd1 vssd1 vccd1 vccd1 _3490_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6671_ net17 _3109_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3883_ _3420_ vssd1 vssd1 vccd1 vccd1 _3421_ sky130_fd_sc_hd__buf_2
X_5622_ _0513_ _0448_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5553_ _1885_ _1886_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__nand2_1
X_4504_ _3406_ _3442_ _0845_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5484_ _1817_ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4435_ _0568_ _0564_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7154_ _0104_ _0265_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_4366_ _0323_ _0708_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _0488_ egd_top.BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _2435_
+ sky130_fd_sc_hd__nand2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _3237_ _3213_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__nand2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7085_ _0035_ _0196_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _1346_ _3349_ _2365_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6938_ _3051_ _3052_ clknet_1_0__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__o21ai_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6869_ clknet_1_0__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__buf_1
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4220_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__clkbuf_4
X_4151_ _0482_ _3282_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__nor2_2
X_4082_ _3226_ _0407_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4984_ _0489_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _1323_
+ sky130_fd_sc_hd__nand2_1
X_3935_ _3217_ _3469_ vssd1 vssd1 vccd1 vccd1 _3473_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6723_ _2810_ _2917_ _2918_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__nand3_1
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6654_ _2803_ _2851_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5605_ _0450_ _0731_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__nand2_1
X_3866_ _3403_ vssd1 vssd1 vccd1 vccd1 _3404_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6585_ _2740_ _2745_ _2784_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3797_ _3334_ vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__buf_2
X_5536_ _3294_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _1870_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5467_ _3195_ _0361_ _3199_ _0364_ _1801_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__a221oi_1
X_4418_ _0503_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _0761_
+ sky130_fd_sc_hd__nand2_1
X_7206_ _0156_ _0317_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dfxtp_2
X_5398_ _1703_ _1733_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__nor2_1
X_7137_ _0087_ _0248_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_4349_ _0678_ _0682_ _0687_ _0691_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__and4_1
X_7068_ _0018_ _0179_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6019_ _3244_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _2349_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__3031_ clknet_0__3031_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3031_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3720_ _3257_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__buf_2
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ _3194_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
X_3582_ _3131_ _3139_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__or2_1
X_6370_ _2628_ _2624_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__and2_1
X_5321_ _1646_ _1649_ _1652_ _1656_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5252_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4203_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__buf_2
Xclkbuf_0__3050_ _3050_ vssd1 vssd1 vccd1 vccd1 clknet_0__3050_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5183_ _3418_ _3401_ _3428_ _3405_ _1519_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__a221oi_1
X_4134_ _0461_ _0464_ _0465_ _0468_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__a221oi_1
X_4065_ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _0877_ _0422_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__or2_1
X_4898_ egd_top.BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__inv_2
X_6706_ _2897_ _2901_ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__nand2_1
X_3918_ _3455_ vssd1 vssd1 vccd1 vccd1 _3456_ sky130_fd_sc_hd__buf_2
X_6637_ _2814_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1
+ vccd1 _2835_ sky130_fd_sc_hd__nand2_1
X_3849_ _3386_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _3387_
+ sky130_fd_sc_hd__nand2_1
X_6568_ _2761_ _2768_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _1210_ _0614_ _1055_ _0618_ _1853_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__a221oi_1
X_6499_ _2713_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5870_ _1589_ _0527_ _0437_ _0530_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4821_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4752_ _3237_ _0801_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3703_ _3240_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__inv_2
X_4683_ _1022_ _0367_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6422_ _2664_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3634_ _3181_ _3166_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__and2_4
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3565_ _3122_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__inv_2
X_6353_ _2616_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6284_ _2569_ _2559_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__and2_1
X_5304_ _3390_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _1640_
+ sky130_fd_sc_hd__nand2_1
X_5235_ _0471_ _3152_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _3335_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _1503_
+ sky130_fd_sc_hd__nand2_1
X_4117_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__clkbuf_4
X_5097_ _1022_ _0422_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__or2_1
X_4048_ _0391_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5999_ _2328_ _2329_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold9 egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _1228_ _1358_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__nor2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6971_ _3023_ vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5922_ egd_top.BitStream_buffer.BS_buffer\[71\] _3378_ _0776_ _3382_ _2252_ vssd1
+ vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5853_ _2183_ _2184_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__nand2_1
X_5784_ _3271_ _3280_ _3285_ _3264_ _2115_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__a221oi_1
X_4804_ _3496_ _3482_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4735_ _1074_ _1075_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4666_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
X_6405_ _2652_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4597_ _0937_ _0603_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__o21ai_1
X_3617_ net5 _3168_ _3159_ vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3548_ _3102_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__inv_2
X_6336_ net13 _0972_ _2469_ vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__mux2_1
X_6267_ net4 _0844_ _2551_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__mux2_1
X_6198_ net8 _3509_ _2479_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__mux2_1
X_5218_ _0695_ _0376_ _3476_ _0379_ _1554_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__a221oi_1
X_5149_ _1359_ _1486_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520_ _0704_ _3502_ _0861_ _3505_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__o22ai_1
X_4451_ _0775_ _0793_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__nand2_1
X_7170_ _0120_ _0281_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3056_ clknet_0__3056_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3056_
+ sky130_fd_sc_hd__clkbuf_16
X_6121_ _2449_ _2450_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__nand2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _0383_ _0382_ _0724_ _0385_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _3366_ _3441_ _2381_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5003_ _0583_ _1073_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6954_ _3054_ _3055_ clknet_1_1__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5905_ _1371_ _3290_ _2235_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__o21ai_1
X_6885_ _3039_ _3040_ clknet_1_1__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5836_ _3205_ _0360_ _3208_ _0363_ _2167_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5767_ _2084_ _2099_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5698_ _1237_ _3501_ _3311_ _3504_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__o22ai_1
X_4718_ egd_top.BitStream_buffer.BS_buffer\[83\] _0494_ _0496_ _1055_ _1058_ vssd1
+ vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4649_ _0679_ _3417_ _0840_ _3421_ _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a221oi_1
X_6319_ _2593_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xsplit1 _3165_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_2
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3951_ _3289_ _3470_ vssd1 vssd1 vccd1 vccd1 _3489_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6670_ _2865_ _2867_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3882_ _3419_ vssd1 vssd1 vccd1 vccd1 _3420_ sky130_fd_sc_hd__clkbuf_2
X_5621_ _0508_ _0442_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__nand2_1
X_5552_ _3389_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _1886_
+ sky130_fd_sc_hd__nand2_1
X_4503_ _3445_ egd_top.BitStream_buffer.BS_buffer\[37\] vssd1 vssd1 vccd1 vccd1 _0845_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5483_ _0456_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _1818_
+ sky130_fd_sc_hd__nand2_1
X_4434_ _0563_ _0551_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4365_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__clkbuf_4
X_7153_ _0103_ _0264_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7084_ _0034_ _0195_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[100\]
+ sky130_fd_sc_hd__dfxtp_1
X_6104_ _2416_ _2433_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__nand2_1
X_4296_ egd_top.BitStream_buffer.BS_buffer\[24\] vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__clkbuf_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _3352_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _2365_
+ sky130_fd_sc_hd__nand2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _3051_ _3052_ clknet_1_0__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6868_ _3027_ vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__buf_4
X_5819_ _3495_ _3512_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__nand2_1
X_6799_ _2971_ _2940_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4150_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__buf_2
X_4081_ egd_top.BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4983_ _1303_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__nand2_1
X_3934_ _3471_ vssd1 vssd1 vccd1 vccd1 _3472_ sky130_fd_sc_hd__buf_2
X_6722_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] _2890_ vssd1 vssd1
+ vccd1 vccd1 _2918_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6653_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__xnor2_1
X_3865_ _3226_ _3398_ vssd1 vssd1 vccd1 vccd1 _3403_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5604_ _0720_ _0426_ _1935_ _1936_ _1937_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__o2111a_1
X_6584_ _2783_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_5_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3796_ _3333_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__clkbuf_2
X_5535_ _0675_ _3253_ _0836_ _3257_ _1868_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5466_ _1157_ _0367_ _1800_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ _0499_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0760_
+ sky130_fd_sc_hd__nand2_1
X_7205_ _0155_ _0316_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dfxtp_2
X_5397_ _1717_ _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__nand2_1
X_7136_ _0086_ _0247_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_4348_ _3453_ _3452_ _3414_ _3456_ _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__a221oi_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7067_ _0017_ _0178_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4279_ _3316_ _0553_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nand2_2
X_6018_ _3236_ _0844_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f__3030_ clknet_0__3030_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3030_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3650_ _3193_ _3166_ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__and2_4
XFILLER_0_43_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3581_ egd_top.BitStream_buffer.pc\[6\] _3107_ _3133_ _3138_ vssd1 vssd1 vccd1 vccd1
+ _3139_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5320_ _3358_ _3452_ _3362_ _3456_ _1655_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5251_ _0448_ _0521_ _0457_ _0525_ _1587_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__a221oi_1
X_4202_ _3260_ _0484_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5182_ _1391_ _3408_ _1518_ _3411_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__o22ai_1
X_4133_ _0472_ _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _3119_ _0407_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6705_ _2898_ _2865_ vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__nand2_1
X_4966_ _0417_ _3171_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__nand2_1
X_4897_ _0844_ _3254_ _0991_ _3258_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__a221oi_1
X_3917_ _3454_ vssd1 vssd1 vccd1 vccd1 _3455_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6636_ _2833_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1
+ vccd1 _2834_ sky130_fd_sc_hd__nand2_1
X_3848_ _3385_ vssd1 vssd1 vccd1 vccd1 _3386_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3779_ _3316_ _3220_ vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6567_ _2767_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5518_ _1729_ _0621_ _1852_ _0624_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__o22ai_1
X_6498_ _2712_ _2689_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__and2_1
X_5449_ _0704_ _3472_ _1781_ _1782_ _1783_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__o2111a_1
X_7119_ _0069_ _0230_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4820_ _3186_ _0348_ _1158_ _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4751_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _3081_ vssd1
+ vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3702_ _3114_ _3230_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__nand2_4
XFILLER_0_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4682_ _0370_ _3174_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6421_ _2663_ _2645_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__and2_1
X_3633_ net16 _3180_ _3159_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3564_ _3119_ _3121_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__nand2_2
X_6352_ _2615_ _2601_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__and2_1
X_6283_ net14 _0675_ _2551_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__mux2_1
X_5303_ _3386_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _1639_
+ sky130_fd_sc_hd__nand2_1
X_5234_ _0741_ _0445_ _0447_ _0894_ _1570_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__a221oi_1
X_5165_ _1491_ _1495_ _1498_ _1501_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__and4_1
Xclkbuf_0__3032_ _3032_ vssd1 vssd1 vccd1 vccd1 clknet_0__3032_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _0442_ _0445_ _0447_ _0448_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5096_ _0417_ _3174_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__nand2_1
X_4047_ _3316_ _0344_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _0567_ _0932_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__nand2_1
X_4949_ _1284_ _1285_ _1286_ _1287_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6619_ _2813_ _2816_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6970_ _3057_ _3058_ clknet_1_0__leaf__3059_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _2250_ _2251_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__nand2_1
X_5852_ _0455_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _2184_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5783_ _1241_ _3290_ _2114_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__o21ai_1
X_4803_ _0855_ _3472_ _1139_ _1140_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__o2111a_1
X_4734_ _0588_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _1075_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4665_ _3468_ _3490_ _0858_ _3493_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6404_ _2651_ _2645_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__and2_1
X_4596_ _0606_ _0597_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__nand2_1
X_3616_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3547_ _3103_ _3104_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__and2b_1
X_6335_ _2604_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6266_ _2557_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
X_6197_ _2509_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
X_5217_ _0700_ _0382_ _0858_ _0385_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o22ai_1
X_5148_ _3212_ _1485_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__nor2_1
X_5079_ _0338_ _3509_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4450_ _0780_ _0785_ _0789_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__and4_1
X_4381_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__inv_2
X_6120_ _0567_ _1073_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__nand2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _3444_ _3372_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__nand2_1
X_5002_ _0615_ _0556_ _0589_ _0560_ _1340_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__a221oi_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6953_ _3054_ _3055_ clknet_1_1__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__o21ai_2
X_5904_ _3294_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _2235_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6884_ _3039_ _3040_ clknet_1_1__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__o21ai_2
X_5835_ _0380_ _0366_ _2166_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5766_ _2088_ _2092_ _2095_ _2098_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__and4_1
X_5697_ _3503_ _3489_ _3500_ _3492_ _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__o221a_1
X_4717_ _1056_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4648_ _0827_ _3424_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__o21ai_1
X_4579_ _0769_ _0528_ _0920_ _0531_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6318_ _2592_ _2580_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__and2_1
X_6249_ _2545_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3950_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _3488_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3881_ _3260_ _3398_ vssd1 vssd1 vccd1 vccd1 _3419_ sky130_fd_sc_hd__and2_1
X_5620_ _0518_ _0493_ _0495_ _0522_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__a221oi_1
X_5551_ _3385_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _1885_
+ sky130_fd_sc_hd__nand2_1
X_4502_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5482_ _0451_ _0413_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__nand2_1
X_4433_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__clkbuf_4
X_4364_ _0705_ _0706_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nor2_1
X_7152_ _0102_ _0263_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_4295_ _3151_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] _3081_ vssd1
+ vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7083_ _0033_ _0194_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[101\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__3038_ clknet_0__3038_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3038_
+ sky130_fd_sc_hd__clkbuf_16
X_6103_ _2420_ _2424_ _2428_ _2432_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__and4_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _0611_ _3325_ _0615_ _3329_ _2363_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__a221oi_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _3051_ _3052_ clknet_1_0__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ _3024_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5818_ _1146_ _3471_ _2147_ _2148_ _2149_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6798_ _2818_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5749_ _0425_ _0543_ _0738_ _0546_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ _0404_ _0409_ _0414_ _0419_ _0423_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4982_ _1307_ _1312_ _1316_ _1320_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3933_ _3234_ _3470_ vssd1 vssd1 vccd1 vccd1 _3471_ sky130_fd_sc_hd__nand2_2
X_6721_ _2890_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1
+ vccd1 vccd1 _2917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3864_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _3402_ sky130_fd_sc_hd__clkbuf_4
X_6652_ _2848_ _2849_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5603_ _0404_ _0438_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6583_ _2778_ _2779_ _2782_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3795_ _3251_ _3121_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__and2_1
X_5534_ _1866_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5465_ _0370_ _3192_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4416_ _0757_ _0486_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__o21ai_1
X_7204_ _0154_ _0315_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7135_ _0085_ _0246_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_2
X_5396_ _1721_ _1725_ _1728_ _1731_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__and4_1
X_4347_ _0688_ _0689_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__nand2_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7066_ _0016_ _0177_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4278_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__inv_2
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6017_ _3150_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] _3161_ vssd1
+ vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__o21ai_1
X_6919_ _3024_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3580_ _3136_ _3137_ _3108_ vssd1 vssd1 vccd1 vccd1 _3138_ sky130_fd_sc_hd__a21oi_1
X_5250_ _0923_ _0528_ _1065_ _0531_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4201_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5181_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__inv_2
X_4132_ _0475_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _0476_
+ sky130_fd_sc_hd__nand2_1
X_4063_ _0406_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__buf_2
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4965_ _0412_ _3163_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__nand2_1
X_6704_ _2897_ _2898_ _2869_ _2867_ _2900_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__a32o_2
X_3916_ _3307_ _3398_ vssd1 vssd1 vccd1 vccd1 _3454_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4896_ _1233_ _1234_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__nand2_1
X_6635_ _2828_ _2829_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__nand2_2
X_3847_ _3384_ vssd1 vssd1 vccd1 vccd1 _3385_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3778_ _3301_ _3231_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__nor2_8
X_6566_ _2765_ _2766_ vssd1 vssd1 vccd1 vccd1 _2767_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5517_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__inv_2
X_6497_ net5 _1073_ _2707_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__mux2_1
X_5448_ _1007_ _3485_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__or2_1
X_5379_ _1589_ _0544_ _0437_ _0547_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_10_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7118_ _0068_ _0229_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_7049_ _3024_ _3027_ clknet_1_0__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4750_ _0951_ _1090_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3701_ _3237_ _3238_ vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4681_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__inv_2
X_6420_ net4 _0452_ _2656_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__mux2_1
X_3632_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__buf_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6351_ net8 _3336_ _2469_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__mux2_1
X_3563_ _3120_ egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\] vssd1
+ vssd1 vccd1 vccd1 _3121_ sky130_fd_sc_hd__and3_2
X_5302_ _3376_ _3361_ _3380_ _3365_ _1637_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__a221oi_1
X_6282_ _2568_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
X_5233_ _1568_ _1569_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__nand2_1
X_5164_ _3439_ _3305_ _0683_ _3310_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__a221oi_1
Xclkbuf_0__3031_ _3031_ vssd1 vssd1 vccd1 vccd1 clknet_0__3031_ sky130_fd_sc_hd__clkbuf_16
X_4115_ _0453_ _0458_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__nand2_1
X_5095_ _0412_ _3168_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__nand2_1
X_4046_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5997_ _0562_ _1073_ vssd1 vssd1 vccd1 vccd1 _2328_ sky130_fd_sc_hd__nand2_1
X_4948_ _0338_ _0865_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__nand2_1
X_4879_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6618_ _2814_ _2815_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6549_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1 vccd1
+ _2750_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__3071_ clknet_0__3071_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3071_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _3389_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _2251_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5851_ _0450_ _0733_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__nand2_1
X_5782_ _3294_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _2114_
+ sky130_fd_sc_hd__nand2_1
X_4802_ _1141_ _3485_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__or2_1
X_4733_ _0583_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _1074_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6403_ net8 _0573_ _2619_ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4664_ _3496_ _3476_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__nand2_1
X_4595_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__inv_2
X_3615_ _3167_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__clkbuf_1
X_3546_ net33 net32 net34 vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__a21o_1
X_6334_ _2603_ _2601_ vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__and2_1
X_6265_ _2556_ _2536_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__and2_1
X_5216_ _3189_ _0361_ _3192_ _0364_ _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6196_ _2492_ _2508_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__and2_1
X_5147_ _1420_ _1483_ _1484_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nand3_2
X_5078_ _0333_ _3275_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__nand2_1
X_4029_ _3168_ _0361_ _3171_ _0364_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4380_ _3171_ _0361_ _3174_ _0364_ _0722_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _3376_ _3416_ _3380_ _3420_ _2379_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__a221oi_1
X_5001_ _1338_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__nand2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6952_ _3054_ _3055_ clknet_1_1__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5903_ _3453_ _3253_ _3414_ _3257_ _2233_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__a221oi_1
X_6883_ _3039_ _3040_ clknet_1_1__leaf__3041_ vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5834_ _0369_ _3202_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5765_ _1192_ _0613_ _0510_ _0617_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5696_ _3495_ _3509_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__nand2_1
X_4716_ _0503_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _1057_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4647_ _3427_ _3372_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4578_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__inv_2
X_6317_ net4 _3362_ _2470_ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__mux2_1
X_3529_ _3089_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__clkbuf_4
X_6248_ _2544_ _2536_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__and2_1
X_6179_ _2497_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3880_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _3418_ sky130_fd_sc_hd__buf_2
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _3322_ _3360_ _3327_ _3364_ _1883_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__a221oi_1
X_5481_ _0365_ _0427_ _1813_ _1814_ _1815_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__o2111a_1
X_4501_ _3428_ _3417_ _0679_ _3421_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4432_ _0767_ _0771_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__and3_1
X_4363_ _3508_ _3512_ _3511_ _3275_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a22o_1
X_7151_ _0101_ _0262_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _3211_ _0637_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__nor2_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7082_ _0032_ _0193_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[102\]
+ sky130_fd_sc_hd__dfxtp_1
X_6102_ _3186_ _0463_ _3189_ _0467_ _2431_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__a221oi_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _1219_ _3122_ _2362_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__o21ai_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6935_ _3051_ _3052_ clknet_1_0__leaf__3053_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__o21ai_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6866_ _3033_ _3034_ clknet_1_1__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__o21ai_2
X_5817_ _0649_ _3484_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__or2_1
X_6797_ _2987_ _2988_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5748_ _0739_ _0520_ _0435_ _0524_ _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_29_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5679_ _3422_ _3407_ _3366_ _3410_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _0733_ _0464_ _3152_ _0468_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6720_ _2914_ _2915_ _2799_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__o21ai_1
X_3932_ _3469_ vssd1 vssd1 vccd1 vccd1 _3470_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6651_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__nand2_1
X_3863_ _3400_ vssd1 vssd1 vccd1 vccd1 _3401_ sky130_fd_sc_hd__buf_2
X_6582_ _2767_ _2780_ _2781_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__a21o_1
X_5602_ _0433_ _3152_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__nand2_1
X_5533_ _3269_ _3395_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__nand2_1
X_3794_ _3122_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _3202_ _0348_ _1797_ _1798_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7203_ _0153_ _0314_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_valid_n
+ sky130_fd_sc_hd__dfxtp_1
X_4415_ _0489_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _0758_
+ sky130_fd_sc_hd__nand2_1
X_5395_ _1073_ _0614_ _1210_ _0618_ _1730_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__a221oi_1
X_7134_ _0084_ _0245_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_4346_ _3463_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0689_
+ sky130_fd_sc_hd__nand2_1
X_7065_ _0015_ _0176_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[80\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4277_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__buf_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6016_ _2226_ _2346_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__nor2_1
X_6918_ _3045_ _3046_ clknet_1_1__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6849_ _3025_ _3028_ clknet_1_0__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _0543_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__buf_2
X_5180_ _1505_ _1509_ _1512_ _1516_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__and4_1
X_4131_ _0474_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4062_ _0405_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4964_ _1294_ _1297_ _1299_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3915_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _3453_ sky130_fd_sc_hd__buf_2
X_6703_ _2899_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4895_ _3270_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _1234_
+ sky130_fd_sc_hd__nand2_1
X_6634_ _2831_ _2813_ _2816_ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__nand3_1
X_3846_ _3316_ _3121_ vssd1 vssd1 vccd1 vccd1 _3384_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3777_ egd_top.BitStream_buffer.BS_buffer\[25\] vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6565_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] vssd1 vssd1 vccd1 vccd1
+ _2766_ sky130_fd_sc_hd__inv_2
X_6496_ _2711_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
X_5516_ _0615_ _0596_ _0589_ _0600_ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__a221oi_1
X_5447_ _3480_ _0865_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__nand2_1
X_5378_ _0457_ _0521_ _0452_ _0525_ _1713_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4329_ _0670_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nand2_1
X_7117_ _0067_ _0228_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_7048_ _3075_ _3076_ clknet_1_0__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3700_ egd_top.BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4680_ _3183_ _0348_ _1019_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__a211oi_1
X_3631_ _3179_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6350_ _2614_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
X_3562_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__inv_2
X_5301_ _0661_ _3368_ _1636_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__o21ai_1
X_6281_ _2567_ _2559_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__and2_1
X_5232_ _0456_ _1039_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__nand2_1
X_5163_ _1371_ _3314_ _1499_ _3318_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_0__3030_ _3030_ vssd1 vssd1 vccd1 vccd1 clknet_0__3030_ sky130_fd_sc_hd__clkbuf_16
X_4114_ _0456_ _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__nand2_1
X_5094_ _1423_ _1426_ _1428_ _1431_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__and4_1
X_4045_ _0388_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__clkbuf_2
X_5996_ _2322_ _2324_ _2326_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__and3_1
X_4947_ _0333_ _3512_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4878_ _0551_ _0596_ _0557_ _0600_ _1217_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6617_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1 vccd1
+ _2815_ sky130_fd_sc_hd__inv_2
X_3829_ _3278_ _3323_ vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6548_ _2747_ _2748_ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6479_ _2702_ _2696_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[3\] sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5850_ _1022_ _0426_ _2179_ _2180_ _2181_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5781_ _3449_ _3253_ _3453_ _3257_ _2112_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4801_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__inv_2
X_4732_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__buf_2
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663_ _0697_ _3472_ _1000_ _1001_ _1003_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__o2111a_1
X_6402_ _2650_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
X_3614_ _3164_ _3166_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__and2_1
X_4594_ _0781_ _0576_ _0932_ _0580_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3545_ _3101_ _3102_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__nor2_1
X_6333_ net14 _0823_ _2470_ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__mux2_1
X_6264_ net5 _0683_ _2551_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5215_ _0873_ _0367_ _1551_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6195_ net9 _0865_ _2479_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__mux2_1
X_5146_ _0633_ _3476_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__nand2_1
X_5077_ _0328_ _3512_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nand2_1
X_4028_ _0365_ _0367_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__o21ai_1
X_5979_ _2308_ _2309_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__3053_ clknet_0__3053_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3053_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _0568_ _0927_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__nand2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6951_ _3054_ _3055_ clknet_1_0__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5902_ _2231_ _2232_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__nand2_1
X_6882_ clknet_1_0__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__buf_1
X_5833_ _0634_ _0347_ _2163_ _2164_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__a211oi_1
X_5764_ _1974_ _0620_ _2096_ _0623_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__o22ai_1
X_5695_ _1007_ _3471_ _2025_ _2026_ _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__o2111a_1
X_4715_ _0499_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _1056_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4646_ _0836_ _3401_ _3449_ _3405_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4577_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _2591_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
X_3528_ _3079_ vssd1 vssd1 vccd1 vccd1 _3089_ sky130_fd_sc_hd__inv_2
X_6247_ net9 _3264_ _2515_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__mux2_1
X_6178_ _2496_ _2492_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__and2_4
X_5129_ _0568_ _0611_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5480_ _0735_ _0439_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__or2_1
X_4500_ _0666_ _3424_ _0841_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__o21ai_1
X_4431_ _0538_ _0537_ _0442_ _0541_ _0773_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _1155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4362_ _3503_ _3502_ _0704_ _3505_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__o22ai_1
X_7150_ _0100_ _0261_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _3212_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__nor2_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7081_ _0031_ _0192_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[103\]
+ sky130_fd_sc_hd__dfxtp_1
X_6101_ _2429_ _2430_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__nand2_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _3334_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _2362_
+ sky130_fd_sc_hd__nand2_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6934_ clknet_1_1__leaf__3031_ vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__buf_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6865_ _3033_ _3034_ clknet_1_1__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__o21ai_2
X_5816_ _3479_ _3275_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6796_ _2966_ _2864_ _2979_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__nand3_1
X_5747_ _1462_ _0527_ _1589_ _0530_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5678_ _2000_ _2003_ _2006_ _2010_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__and4_1
X_4629_ _0657_ _3326_ _0818_ _3330_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4980_ _1317_ _1318_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__nand2_1
X_3931_ _3120_ _3396_ _3218_ vssd1 vssd1 vccd1 vccd1 _3469_ sky130_fd_sc_hd__and3_2
XFILLER_0_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6650_ _2847_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3862_ _3399_ vssd1 vssd1 vccd1 vccd1 _3400_ sky130_fd_sc_hd__clkbuf_2
X_6581_ _2772_ _3150_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__nand2_1
X_5601_ _0429_ _0418_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__nand2_1
X_5532_ _3262_ _3402_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__nand2_1
X_3793_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5463_ _0354_ egd_top.BitStream_buffer.BS_buffer\[127\] _0356_ egd_top.BitStream_buffer.BS_buffer\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4414_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__inv_2
X_5394_ _1605_ _0621_ _1729_ _0624_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__o22ai_1
X_7202_ _0152_ _0313_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7133_ _0083_ _0244_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_4345_ _3459_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _0688_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7064_ _0014_ _0175_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[81\]
+ sky130_fd_sc_hd__dfxtp_1
X_4276_ _3312_ _0553_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__nand2_2
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6015_ _3149_ _2345_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6917_ _3045_ _3046_ clknet_1_1__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__o21ai_2
X_6848_ _3025_ _3028_ clknet_1_1__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6779_ _2971_ vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4130_ _0473_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__clkbuf_2
X_4061_ egd_top.BitStream_buffer.pc\[4\] _3120_ _3218_ vssd1 vssd1 vccd1 vccd1 _0405_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ _3202_ _0390_ _3205_ _0393_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6702_ _2743_ net18 _2744_ _3110_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3914_ _3451_ vssd1 vssd1 vccd1 vccd1 _3452_ sky130_fd_sc_hd__buf_2
X_4894_ _3263_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _1233_
+ sky130_fd_sc_hd__nand2_1
X_6633_ _2827_ _2830_ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3845_ _3382_ vssd1 vssd1 vccd1 vccd1 _3383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3776_ _3313_ vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__buf_2
X_6564_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] _2764_ vssd1 vssd1
+ vccd1 vccd1 _2765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6495_ _2710_ _2689_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__and2_1
X_5515_ _0622_ _0603_ _1849_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ _3475_ _3512_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__nand2_1
X_5377_ _1065_ _0528_ _1202_ _0531_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__o22ai_1
X_4328_ _3390_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0671_
+ sky130_fd_sc_hd__nand2_1
X_7116_ _0066_ _0227_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_7047_ _3075_ _3076_ clknet_1_0__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__o21ai_2
X_4259_ _0602_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__buf_2
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3630_ _3178_ _3166_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__and2_1
X_3561_ _3118_ vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__buf_6
X_5300_ _3371_ _0972_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__nand2_1
X_6280_ net15 _3402_ _2551_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5231_ _0451_ _0461_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__nand2_1
X_5162_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__inv_2
X_4113_ egd_top.BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__clkbuf_4
X_5093_ _3205_ _0390_ _3208_ _0393_ _1430_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__a221oi_1
X_4044_ _3312_ _0344_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5995_ _0465_ _0536_ _0413_ _0540_ _2325_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__a221oi_1
X_4946_ _0328_ _3509_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4877_ _1215_ _0603_ _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6616_ _2797_ _2809_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__nor2_4
X_3828_ egd_top.BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _3366_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6547_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1 vccd1
+ _2748_ sky130_fd_sc_hd__inv_2
X_3759_ _3295_ _3296_ vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__nand2_1
X_6478_ _2697_ _2698_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__nand2_2
X_5429_ _1762_ _1763_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _3480_ _0339_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5780_ _2110_ _2111_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4731_ _0927_ _0556_ _0611_ _0560_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__a221oi_1
X_4662_ _1002_ _3485_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6401_ _2649_ _2645_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__and2_1
X_3613_ _3165_ vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__buf_6
X_4593_ _0933_ _0934_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nand2_1
X_3544_ net33 net32 vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6332_ _2602_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
X_6263_ _2555_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5214_ _0370_ _3186_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6194_ _2507_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__clkbuf_1
X_5145_ _1450_ _1482_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5076_ _0323_ _3287_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__nand2_1
X_4027_ _0370_ _3163_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5978_ _0474_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _2309_
+ sky130_fd_sc_hd__nand2_1
X_4929_ _0837_ _3442_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6950_ _3054_ _3055_ clknet_1_0__leaf__3056_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__o21ai_2
X_5901_ _3269_ _0836_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6881_ _3027_ vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__buf_4
X_5832_ _0353_ _0947_ _0355_ _3497_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5763_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4714_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__clkbuf_4
X_5694_ _3288_ _3484_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__or2_1
X_4645_ _0837_ _3408_ _0985_ _3411_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4576_ _0910_ _0914_ _0915_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__and4b_1
X_3527_ net38 net37 vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__nand2_1
X_6315_ _2590_ _2580_ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__and2_1
X_6246_ _2543_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
X_6177_ net15 _3482_ _2480_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__mux2_1
X_5128_ _0563_ _0615_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _3445_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _1397_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4430_ _0545_ _0544_ _0772_ _0547_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__o22ai_1
XANTENNA_2 _1419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__3035_ clknet_0__3035_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3035_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6100_ _0474_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _2430_
+ sky130_fd_sc_hd__nand2_1
X_4361_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7080_ _0030_ _0191_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[104\]
+ sky130_fd_sc_hd__dfxtp_1
X_4292_ _0343_ _0629_ _0635_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__nand3_2
X_6031_ _2351_ _2355_ _2358_ _2360_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__and4_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6933_ _3027_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__buf_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6864_ _3033_ _3034_ clknet_1_1__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__o21ai_2
X_5815_ _3474_ _0648_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6795_ _2958_ _2986_ _2865_ vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5746_ _2072_ _2076_ _2077_ _2078_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__and4b_1
X_5677_ _0564_ _3378_ _0551_ _3382_ _2009_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__a221oi_1
X_4628_ _0937_ _3332_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__o21ai_1
X_4559_ _0457_ _0445_ _0447_ _0452_ _0900_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a221oi_1
X_6229_ _2513_ _2531_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__and2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3930_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _3468_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3861_ _3217_ _3398_ vssd1 vssd1 vccd1 vccd1 _3399_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6580_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2780_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3792_ _3329_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__buf_2
X_5600_ _1157_ _0408_ _1931_ _1932_ _1933_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__o2111a_1
X_5531_ _3432_ _3222_ _3439_ _3228_ _1864_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7201_ _0151_ _0312_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[113\]
+ sky130_fd_sc_hd__dfxtp_1
X_5462_ _0724_ _0351_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5393_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__inv_2
X_4413_ _0730_ _0755_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7132_ _0082_ _0243_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_4344_ _3439_ _3435_ _3438_ _0683_ _0686_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__a221oi_1
X_7063_ _0013_ _0174_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[82\]
+ sky130_fd_sc_hd__dfxtp_1
X_4275_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__inv_2
X_6014_ _2283_ _2343_ _2344_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__nand3_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6916_ _3045_ _3046_ clknet_1_1__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6847_ _3025_ _3028_ clknet_1_1__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6778_ _2814_ _2754_ _2758_ vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5729_ _0455_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _2062_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4060_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__inv_2
X_4962_ _1026_ _0396_ _1300_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__o21ai_1
X_4893_ _3306_ _3223_ _3271_ _3229_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__a221oi_1
X_6701_ _2895_ _2861_ _2860_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__nand3_1
X_3913_ _3450_ vssd1 vssd1 vccd1 vccd1 _3451_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6632_ _2828_ _2746_ _2829_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__nand3_1
X_3844_ _3381_ vssd1 vssd1 vccd1 vccd1 _3382_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3775_ _3312_ _3220_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__nand2_2
X_6563_ _2762_ _2763_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6494_ net6 _0932_ _2707_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5514_ _0606_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _1849_
+ sky130_fd_sc_hd__nand2_1
X_5445_ _1769_ _1772_ _1775_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5376_ _1705_ _1709_ _1710_ _1711_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__and4b_1
X_7115_ _0065_ _0226_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_4327_ _3386_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _0670_
+ sky130_fd_sc_hd__nand2_1
X_7046_ _3075_ _3076_ clknet_1_0__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__o21ai_2
X_4258_ _3278_ _0553_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__nand2_2
X_4189_ _0518_ _0521_ _0522_ _0525_ _0532_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3560_ _3117_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1
+ vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__and3_1
X_5230_ _0735_ _0427_ _1564_ _1565_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__o2111a_1
X_5161_ _3224_ _3281_ _3286_ _0639_ _1497_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__buf_2
X_5092_ _3491_ _0396_ _1429_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__o21ai_1
X_4043_ _3205_ _0376_ _3208_ _0379_ _0386_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__a221oi_1
X_5994_ _0892_ _0543_ _1037_ _0546_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__o22ai_1
X_4945_ _0323_ _3275_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4876_ _0606_ _0564_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6615_ _2797_ _2809_ _2748_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__o21ai_1
X_3827_ _3364_ vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__buf_2
X_3758_ egd_top.BitStream_buffer.BS_buffer\[19\] vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__clkbuf_4
X_6546_ _2746_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1
+ vccd1 _2747_ sky130_fd_sc_hd__nand2_1
X_3689_ _3226_ _3220_ vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__and2_1
X_6477_ _3396_ _3090_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__nor2_1
X_5428_ _3390_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _1763_
+ sky130_fd_sc_hd__nand2_1
X_5359_ _0456_ _0461_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__nand2_1
X_7029_ _3072_ _3073_ clknet_1_1__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4730_ _1069_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4661_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6400_ net9 _0584_ _2619_ vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__mux2_1
X_3612_ _3079_ vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__buf_8
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4592_ _0588_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _0934_
+ sky130_fd_sc_hd__nand2_1
X_6331_ _2600_ _2601_ vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__and2_1
X_3543_ net34 vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__inv_2
X_6262_ _2554_ _2536_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5213_ _3195_ _0348_ _1548_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__a211oi_1
X_6193_ _2506_ _2492_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__and2_4
X_5144_ _1465_ _1481_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5075_ _1411_ _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4026_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__buf_2
X_5977_ _0470_ _3180_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__nand2_1
X_4928_ _3445_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _1267_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4859_ _1191_ _1196_ _1197_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__and4b_1
X_6529_ _2733_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5900_ _3262_ _3449_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6880_ _3024_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__buf_4
X_5831_ _3491_ _0350_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__nor2_1
X_5762_ _0584_ _0595_ _0573_ _0599_ _2094_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4713_ _0526_ _0486_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5693_ _3479_ _3512_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4644_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4575_ _0514_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3526_ _3082_ _3083_ _3085_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__a21o_1
X_6314_ net5 _3358_ _2470_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__mux2_1
X_6245_ _2542_ _2536_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__and2_1
X_6176_ _2495_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
X_5127_ _1459_ _1461_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__and3_1
X_5058_ _3358_ _3417_ _3362_ _3421_ _1395_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__a221oi_1
X_4009_ _3217_ _0345_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_3 _2282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4360_ _0700_ _3490_ _3488_ _3493_ _0702_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__o221a_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _0633_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__nand2_1
X_6030_ _0675_ _3304_ _0836_ _3309_ _2359_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__a221oi_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6932_ _3024_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__buf_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6863_ _3033_ _3034_ clknet_1_0__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__o21ai_2
X_5814_ _2135_ _2138_ _2141_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6794_ _2978_ _2861_ _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__nand3_1
XFILLER_0_29_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5745_ _0513_ _0457_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__nand2_1
X_5676_ _2007_ _2008_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4627_ _3335_ _0607_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4558_ _0898_ _0899_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__nand2_1
X_4489_ _3386_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _0831_
+ sky130_fd_sc_hd__nand2_1
X_6228_ net15 _3224_ _2516_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__mux2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _2483_ _3197_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__and2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3860_ _3397_ vssd1 vssd1 vccd1 vccd1 _3398_ sky130_fd_sc_hd__clkbuf_4
X_3791_ _3328_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__clkbuf_2
X_5530_ _1862_ _1863_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5461_ _1752_ _1766_ _1780_ _1795_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__and4_1
X_4412_ _0737_ _0745_ _0750_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__and4_1
X_7200_ _0150_ _0311_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[114\]
+ sky130_fd_sc_hd__dfxtp_1
X_5392_ _0611_ _0596_ _0615_ _0600_ _1727_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4343_ _0684_ _3442_ _0685_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__o21ai_1
X_7131_ _0081_ _0242_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_7062_ _0012_ _0173_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[83\]
+ sky130_fd_sc_hd__dfxtp_1
X_4274_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__buf_2
X_6013_ _0632_ _0865_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__nand2_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6915_ _3045_ _3046_ clknet_1_1__leaf__3047_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6846_ _3025_ _3028_ clknet_1_1__leaf__3032_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__o21ai_2
X_6777_ _2903_ _2969_ _2941_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__nand3_1
X_3989_ _0332_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5728_ _0450_ _0418_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5659_ _3294_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _1992_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ _0399_ _3208_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__nand2_1
X_4892_ _1229_ _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6700_ _2896_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3912_ _3302_ _3397_ vssd1 vssd1 vccd1 vccd1 _3450_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6631_ _2797_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__inv_2
X_3843_ _3307_ _3323_ vssd1 vssd1 vccd1 vccd1 _3381_ sky130_fd_sc_hd__and2_1
X_3774_ _3301_ _3240_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__nor2_8
X_6562_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] vssd1 vssd1 vccd1 vccd1
+ _2763_ sky130_fd_sc_hd__inv_4
X_5513_ _0515_ _0576_ _0765_ _0580_ _1847_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__a221oi_1
X_6493_ _2709_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5444_ _3362_ _3452_ _3340_ _3456_ _1778_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5375_ _0514_ _0538_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__nand2_1
X_7114_ _0064_ _0225_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ _3362_ _3361_ _3340_ _3365_ _0668_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__a221oi_1
X_7045_ _3075_ _3076_ clknet_1_0__leaf__3077_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__o21ai_2
X_4257_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__inv_2
X_4188_ _0526_ _0528_ _0529_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6829_ _3013_ _3019_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__3068_ clknet_0__3068_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__3068_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5160_ _3315_ _3291_ _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__o21ai_1
X_4111_ _0454_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__clkbuf_2
X_5091_ _0399_ _0634_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__nand2_1
X_4042_ _0380_ _0382_ _0383_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__o22ai_1
X_5993_ _0741_ _0520_ _0894_ _0524_ _2323_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__a221oi_1
X_4944_ _1281_ _1282_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4875_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6614_ _2807_ _2808_ _2811_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__a21oi_1
X_3826_ _3363_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__clkbuf_2
X_3757_ _3294_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6545_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1 vccd1
+ _2746_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3688_ _3225_ vssd1 vssd1 vccd1 vccd1 _3226_ sky130_fd_sc_hd__buf_4
X_6476_ egd_top.BitStream_buffer.pc_previous\[4\] _2699_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[4\]
+ sky130_fd_sc_hd__xor2_2
X_5427_ _3386_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _1762_
+ sky130_fd_sc_hd__nand2_1
X_5358_ _0451_ _0465_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__nand2_1
X_4309_ _3287_ _3281_ _3286_ _0648_ _0651_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__a221oi_1
X_5289_ _0639_ _3281_ _3286_ _0801_ _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__a221oi_1
X_7028_ _3072_ _3073_ clknet_1_0__leaf__3074_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_65_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4660_ _3480_ _3482_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611_ net6 _3163_ _3159_ vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__mux2_1
X_4591_ _0583_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _0933_
+ sky130_fd_sc_hd__nand2_1
X_6330_ net39 vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__clkbuf_2
X_3542_ _3100_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__inv_2
X_6261_ net6 _3439_ _2551_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__mux2_1
X_5212_ _0354_ _3202_ _0356_ _3205_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__a22o_1
X_6192_ net10 _0708_ _2479_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5143_ _1469_ _1473_ _1477_ _1480_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__and4_1
X_5074_ _3508_ _3246_ _3511_ _3238_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5976_ _0731_ _0444_ _0446_ _0418_ _2306_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__a221oi_1
X_4927_ _3372_ _3417_ _3358_ _3421_ _1265_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__a221oi_1
X_4858_ _0514_ _0522_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__nand2_1
X_3809_ _3346_ vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__buf_2
XFILLER_0_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4789_ _0840_ _3417_ _3372_ _3421_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__a221oi_1
X_6528_ _2732_ _3080_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6459_ _2688_ _2689_ vssd1 vssd1 vccd1 vccd1 _2690_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__3050_ clknet_0__3050_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__3050_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5830_ _2119_ _2133_ _2146_ _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__and4_1
X_5761_ _0941_ _0602_ _2093_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__o21ai_1
X_4712_ _0489_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _1053_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5692_ _3474_ _3287_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4643_ _0970_ _0975_ _0979_ _0983_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4574_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__clkbuf_4
X_3525_ _3086_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
X_6313_ _2589_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
X_6244_ net10 _3271_ _2515_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6175_ _2492_ _2494_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__and2_1
X_5126_ _0746_ _0537_ _0739_ _0541_ _1463_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__a221oi_1
X_5057_ _1252_ _3424_ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__o21ai_1
X_4008_ _0349_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5959_ _0855_ _0381_ _1002_ _0384_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _3026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__clkbuf_4
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6931_ _3048_ _3049_ clknet_1_1__leaf__3050_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__o21ai_2
X_6862_ _3033_ _3034_ clknet_1_1__leaf__3035_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5813_ _3354_ _3451_ _0662_ _3455_ _2144_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__a221oi_1
X_6793_ _2945_ _2953_ vssd1 vssd1 vccd1 vccd1 _2985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5744_ _0508_ _0448_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5675_ _3389_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _2008_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4626_ _0955_ _0959_ _0963_ _0966_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__and4_1
XFILLER_0_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4557_ _0456_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _0899_
+ sky130_fd_sc_hd__nand2_1
X_4488_ _3340_ _3361_ _3344_ _3365_ _0829_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__a221oi_1
X_6227_ _2530_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ net6 _0796_ _2480_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__mux2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _1445_ _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__nand2_1
X_6089_ _0394_ _0421_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 la_data_out_15_8[6] sky130_fd_sc_hd__buf_12
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _3260_ _3323_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5460_ _1784_ _1786_ _1789_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4411_ _0465_ _0464_ _0413_ _0468_ _0753_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5391_ _0619_ _0603_ _1726_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4342_ _3445_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _0685_
+ sky130_fd_sc_hd__nand2_1
X_7130_ _0080_ _0241_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7061_ _0011_ _0172_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[84\]
+ sky130_fd_sc_hd__dfxtp_2
X_4273_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__clkbuf_2
X_6012_ _2313_ _2342_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__nor2_1
.ends

