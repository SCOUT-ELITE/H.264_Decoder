// This is the unpowered netlist.
module egd_top_wrapper (la_data_in_65,
    wb_clk_i,
    la_data_in_47_32,
    la_data_in_49_48,
    la_data_out_15_8,
    la_data_out_18_16,
    la_data_out_22_19);
 input la_data_in_65;
 input wb_clk_i;
 input [15:0] la_data_in_47_32;
 input [1:0] la_data_in_49_48;
 output [7:0] la_data_out_15_8;
 output [2:0] la_data_out_18_16;
 output [3:0] la_data_out_22_19;

 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire clknet_0__2717_;
 wire clknet_0__2718_;
 wire clknet_0__2719_;
 wire clknet_0__2720_;
 wire clknet_0__2721_;
 wire clknet_0__2722_;
 wire clknet_0__2723_;
 wire clknet_0__2724_;
 wire clknet_0__2725_;
 wire clknet_0__2726_;
 wire clknet_0__2727_;
 wire clknet_0__2728_;
 wire clknet_0__2729_;
 wire clknet_0__2730_;
 wire clknet_0__2731_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf__2717_;
 wire clknet_1_0__leaf__2718_;
 wire clknet_1_0__leaf__2719_;
 wire clknet_1_0__leaf__2720_;
 wire clknet_1_0__leaf__2721_;
 wire clknet_1_0__leaf__2722_;
 wire clknet_1_0__leaf__2723_;
 wire clknet_1_0__leaf__2724_;
 wire clknet_1_0__leaf__2725_;
 wire clknet_1_0__leaf__2726_;
 wire clknet_1_0__leaf__2727_;
 wire clknet_1_0__leaf__2728_;
 wire clknet_1_0__leaf__2729_;
 wire clknet_1_0__leaf__2730_;
 wire clknet_1_0__leaf__2731_;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf__2717_;
 wire clknet_1_1__leaf__2718_;
 wire clknet_1_1__leaf__2719_;
 wire clknet_1_1__leaf__2720_;
 wire clknet_1_1__leaf__2721_;
 wire clknet_1_1__leaf__2722_;
 wire clknet_1_1__leaf__2723_;
 wire clknet_1_1__leaf__2724_;
 wire clknet_1_1__leaf__2725_;
 wire clknet_1_1__leaf__2726_;
 wire clknet_1_1__leaf__2727_;
 wire clknet_1_1__leaf__2728_;
 wire clknet_1_1__leaf__2729_;
 wire clknet_1_1__leaf__2730_;
 wire clknet_1_1__leaf__2731_;
 wire clknet_1_1__leaf_wb_clk_i;
 wire \egd_top.BitStream_buffer.BS_buffer[0] ;
 wire \egd_top.BitStream_buffer.BS_buffer[100] ;
 wire \egd_top.BitStream_buffer.BS_buffer[101] ;
 wire \egd_top.BitStream_buffer.BS_buffer[102] ;
 wire \egd_top.BitStream_buffer.BS_buffer[103] ;
 wire \egd_top.BitStream_buffer.BS_buffer[104] ;
 wire \egd_top.BitStream_buffer.BS_buffer[105] ;
 wire \egd_top.BitStream_buffer.BS_buffer[106] ;
 wire \egd_top.BitStream_buffer.BS_buffer[107] ;
 wire \egd_top.BitStream_buffer.BS_buffer[108] ;
 wire \egd_top.BitStream_buffer.BS_buffer[109] ;
 wire \egd_top.BitStream_buffer.BS_buffer[10] ;
 wire \egd_top.BitStream_buffer.BS_buffer[110] ;
 wire \egd_top.BitStream_buffer.BS_buffer[111] ;
 wire \egd_top.BitStream_buffer.BS_buffer[112] ;
 wire \egd_top.BitStream_buffer.BS_buffer[113] ;
 wire \egd_top.BitStream_buffer.BS_buffer[114] ;
 wire \egd_top.BitStream_buffer.BS_buffer[115] ;
 wire \egd_top.BitStream_buffer.BS_buffer[116] ;
 wire \egd_top.BitStream_buffer.BS_buffer[117] ;
 wire \egd_top.BitStream_buffer.BS_buffer[118] ;
 wire \egd_top.BitStream_buffer.BS_buffer[119] ;
 wire \egd_top.BitStream_buffer.BS_buffer[11] ;
 wire \egd_top.BitStream_buffer.BS_buffer[120] ;
 wire \egd_top.BitStream_buffer.BS_buffer[121] ;
 wire \egd_top.BitStream_buffer.BS_buffer[122] ;
 wire \egd_top.BitStream_buffer.BS_buffer[123] ;
 wire \egd_top.BitStream_buffer.BS_buffer[124] ;
 wire \egd_top.BitStream_buffer.BS_buffer[125] ;
 wire \egd_top.BitStream_buffer.BS_buffer[126] ;
 wire \egd_top.BitStream_buffer.BS_buffer[127] ;
 wire \egd_top.BitStream_buffer.BS_buffer[12] ;
 wire \egd_top.BitStream_buffer.BS_buffer[13] ;
 wire \egd_top.BitStream_buffer.BS_buffer[14] ;
 wire \egd_top.BitStream_buffer.BS_buffer[15] ;
 wire \egd_top.BitStream_buffer.BS_buffer[16] ;
 wire \egd_top.BitStream_buffer.BS_buffer[17] ;
 wire \egd_top.BitStream_buffer.BS_buffer[18] ;
 wire \egd_top.BitStream_buffer.BS_buffer[19] ;
 wire \egd_top.BitStream_buffer.BS_buffer[1] ;
 wire \egd_top.BitStream_buffer.BS_buffer[20] ;
 wire \egd_top.BitStream_buffer.BS_buffer[21] ;
 wire \egd_top.BitStream_buffer.BS_buffer[22] ;
 wire \egd_top.BitStream_buffer.BS_buffer[23] ;
 wire \egd_top.BitStream_buffer.BS_buffer[24] ;
 wire \egd_top.BitStream_buffer.BS_buffer[25] ;
 wire \egd_top.BitStream_buffer.BS_buffer[26] ;
 wire \egd_top.BitStream_buffer.BS_buffer[27] ;
 wire \egd_top.BitStream_buffer.BS_buffer[28] ;
 wire \egd_top.BitStream_buffer.BS_buffer[29] ;
 wire \egd_top.BitStream_buffer.BS_buffer[2] ;
 wire \egd_top.BitStream_buffer.BS_buffer[30] ;
 wire \egd_top.BitStream_buffer.BS_buffer[31] ;
 wire \egd_top.BitStream_buffer.BS_buffer[32] ;
 wire \egd_top.BitStream_buffer.BS_buffer[33] ;
 wire \egd_top.BitStream_buffer.BS_buffer[34] ;
 wire \egd_top.BitStream_buffer.BS_buffer[35] ;
 wire \egd_top.BitStream_buffer.BS_buffer[36] ;
 wire \egd_top.BitStream_buffer.BS_buffer[37] ;
 wire \egd_top.BitStream_buffer.BS_buffer[38] ;
 wire \egd_top.BitStream_buffer.BS_buffer[39] ;
 wire \egd_top.BitStream_buffer.BS_buffer[3] ;
 wire \egd_top.BitStream_buffer.BS_buffer[40] ;
 wire \egd_top.BitStream_buffer.BS_buffer[41] ;
 wire \egd_top.BitStream_buffer.BS_buffer[42] ;
 wire \egd_top.BitStream_buffer.BS_buffer[43] ;
 wire \egd_top.BitStream_buffer.BS_buffer[44] ;
 wire \egd_top.BitStream_buffer.BS_buffer[45] ;
 wire \egd_top.BitStream_buffer.BS_buffer[46] ;
 wire \egd_top.BitStream_buffer.BS_buffer[47] ;
 wire \egd_top.BitStream_buffer.BS_buffer[48] ;
 wire \egd_top.BitStream_buffer.BS_buffer[49] ;
 wire \egd_top.BitStream_buffer.BS_buffer[4] ;
 wire \egd_top.BitStream_buffer.BS_buffer[50] ;
 wire \egd_top.BitStream_buffer.BS_buffer[51] ;
 wire \egd_top.BitStream_buffer.BS_buffer[52] ;
 wire \egd_top.BitStream_buffer.BS_buffer[53] ;
 wire \egd_top.BitStream_buffer.BS_buffer[54] ;
 wire \egd_top.BitStream_buffer.BS_buffer[55] ;
 wire \egd_top.BitStream_buffer.BS_buffer[56] ;
 wire \egd_top.BitStream_buffer.BS_buffer[57] ;
 wire \egd_top.BitStream_buffer.BS_buffer[58] ;
 wire \egd_top.BitStream_buffer.BS_buffer[59] ;
 wire \egd_top.BitStream_buffer.BS_buffer[5] ;
 wire \egd_top.BitStream_buffer.BS_buffer[60] ;
 wire \egd_top.BitStream_buffer.BS_buffer[61] ;
 wire \egd_top.BitStream_buffer.BS_buffer[62] ;
 wire \egd_top.BitStream_buffer.BS_buffer[63] ;
 wire \egd_top.BitStream_buffer.BS_buffer[64] ;
 wire \egd_top.BitStream_buffer.BS_buffer[65] ;
 wire \egd_top.BitStream_buffer.BS_buffer[66] ;
 wire \egd_top.BitStream_buffer.BS_buffer[67] ;
 wire \egd_top.BitStream_buffer.BS_buffer[68] ;
 wire \egd_top.BitStream_buffer.BS_buffer[69] ;
 wire \egd_top.BitStream_buffer.BS_buffer[6] ;
 wire \egd_top.BitStream_buffer.BS_buffer[70] ;
 wire \egd_top.BitStream_buffer.BS_buffer[71] ;
 wire \egd_top.BitStream_buffer.BS_buffer[72] ;
 wire \egd_top.BitStream_buffer.BS_buffer[73] ;
 wire \egd_top.BitStream_buffer.BS_buffer[74] ;
 wire \egd_top.BitStream_buffer.BS_buffer[75] ;
 wire \egd_top.BitStream_buffer.BS_buffer[76] ;
 wire \egd_top.BitStream_buffer.BS_buffer[77] ;
 wire \egd_top.BitStream_buffer.BS_buffer[78] ;
 wire \egd_top.BitStream_buffer.BS_buffer[79] ;
 wire \egd_top.BitStream_buffer.BS_buffer[7] ;
 wire \egd_top.BitStream_buffer.BS_buffer[80] ;
 wire \egd_top.BitStream_buffer.BS_buffer[81] ;
 wire \egd_top.BitStream_buffer.BS_buffer[82] ;
 wire \egd_top.BitStream_buffer.BS_buffer[83] ;
 wire \egd_top.BitStream_buffer.BS_buffer[84] ;
 wire \egd_top.BitStream_buffer.BS_buffer[85] ;
 wire \egd_top.BitStream_buffer.BS_buffer[86] ;
 wire \egd_top.BitStream_buffer.BS_buffer[87] ;
 wire \egd_top.BitStream_buffer.BS_buffer[88] ;
 wire \egd_top.BitStream_buffer.BS_buffer[89] ;
 wire \egd_top.BitStream_buffer.BS_buffer[8] ;
 wire \egd_top.BitStream_buffer.BS_buffer[90] ;
 wire \egd_top.BitStream_buffer.BS_buffer[91] ;
 wire \egd_top.BitStream_buffer.BS_buffer[92] ;
 wire \egd_top.BitStream_buffer.BS_buffer[93] ;
 wire \egd_top.BitStream_buffer.BS_buffer[94] ;
 wire \egd_top.BitStream_buffer.BS_buffer[95] ;
 wire \egd_top.BitStream_buffer.BS_buffer[96] ;
 wire \egd_top.BitStream_buffer.BS_buffer[97] ;
 wire \egd_top.BitStream_buffer.BS_buffer[98] ;
 wire \egd_top.BitStream_buffer.BS_buffer[99] ;
 wire \egd_top.BitStream_buffer.BS_buffer[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[10] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[11] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[12] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[13] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[14] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[15] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[1] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[2] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[3] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[4] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[5] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[6] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[7] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[8] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_output[9] ;
 wire \egd_top.BitStream_buffer.BitStream_buffer_valid_n ;
 wire \egd_top.BitStream_buffer.buffer_index[4] ;
 wire \egd_top.BitStream_buffer.buffer_index[5] ;
 wire \egd_top.BitStream_buffer.buffer_index[6] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[1] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[2] ;
 wire \egd_top.BitStream_buffer.exp_golomb_len[3] ;
 wire \egd_top.BitStream_buffer.pc[0] ;
 wire \egd_top.BitStream_buffer.pc[1] ;
 wire \egd_top.BitStream_buffer.pc[2] ;
 wire \egd_top.BitStream_buffer.pc[3] ;
 wire \egd_top.BitStream_buffer.pc[4] ;
 wire \egd_top.BitStream_buffer.pc[5] ;
 wire \egd_top.BitStream_buffer.pc[6] ;
 wire \egd_top.BitStream_buffer.pc_previous[0] ;
 wire \egd_top.BitStream_buffer.pc_previous[1] ;
 wire \egd_top.BitStream_buffer.pc_previous[2] ;
 wire \egd_top.BitStream_buffer.pc_previous[3] ;
 wire \egd_top.BitStream_buffer.pc_previous[4] ;
 wire \egd_top.BitStream_buffer.pc_previous[5] ;
 wire \egd_top.BitStream_buffer.pc_previous[6] ;
 wire \egd_top.BitStream_buffer.pc_reg[0] ;
 wire \egd_top.BitStream_buffer.pc_reg[1] ;
 wire \egd_top.BitStream_buffer.pc_reg[2] ;
 wire \egd_top.BitStream_buffer.pc_reg[3] ;
 wire \egd_top.BitStream_buffer.pc_reg[4] ;
 wire \egd_top.BitStream_buffer.pc_reg[5] ;
 wire \egd_top.BitStream_buffer.pc_reg[6] ;
 wire \egd_top.exp_golomb_decoding.te_range[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_1206_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_1495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_1767_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_2064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_2160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_2162_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_2276_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_2771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_2864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_2979_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_3031_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_3078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_3078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_3101_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_0583_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_2816_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_2895_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0505_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0757_));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_88 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3158_ (.A(net33),
    .Y(_2732_));
 sky130_fd_sc_hd__nand2_1 _3159_ (.A(net32),
    .B(net31),
    .Y(_2733_));
 sky130_fd_sc_hd__inv_2 _3160_ (.A(net222),
    .Y(_2734_));
 sky130_fd_sc_hd__o21ai_1 _3161_ (.A1(_2732_),
    .A2(_2733_),
    .B1(_2734_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_1 _3162_ (.A(net33),
    .B(net32),
    .Y(_2735_));
 sky130_fd_sc_hd__nor2_1 _3163_ (.A(_2734_),
    .B(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__inv_2 _3164_ (.A(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__a21o_1 _3165_ (.A1(_2732_),
    .A2(_2733_),
    .B1(_0328_),
    .X(_2738_));
 sky130_fd_sc_hd__o21ai_1 _3166_ (.A1(_2732_),
    .A2(_2737_),
    .B1(_2738_),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _3167_ (.A(net31),
    .Y(_2739_));
 sky130_fd_sc_hd__nor2_1 _3168_ (.A(_2739_),
    .B(_2736_),
    .Y(_2740_));
 sky130_fd_sc_hd__o22a_1 _3169_ (.A1(_2733_),
    .A2(_2736_),
    .B1(net32),
    .B2(_2740_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_1 _3170_ (.A(net31),
    .B(_2737_),
    .Y(_2741_));
 sky130_fd_sc_hd__nor2_1 _3171_ (.A(_2740_),
    .B(_2741_),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _3172_ (.A(net30),
    .Y(_2742_));
 sky130_fd_sc_hd__inv_2 _3173_ (.A(net28),
    .Y(_2743_));
 sky130_fd_sc_hd__inv_2 _3174_ (.A(net29),
    .Y(_2744_));
 sky130_fd_sc_hd__nand2_1 _3175_ (.A(_2742_),
    .B(_2744_),
    .Y(_2745_));
 sky130_fd_sc_hd__nand2_1 _3176_ (.A(_2743_),
    .B(net29),
    .Y(_2746_));
 sky130_fd_sc_hd__o211a_1 _3177_ (.A1(_2742_),
    .A2(_2743_),
    .B1(_2745_),
    .C1(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__nand2_1 _3178_ (.A(_2744_),
    .B(net28),
    .Y(_2748_));
 sky130_fd_sc_hd__nand2_1 _3179_ (.A(net30),
    .B(net29),
    .Y(_2749_));
 sky130_fd_sc_hd__nor2_1 _3180_ (.A(net28),
    .B(_2745_),
    .Y(_2750_));
 sky130_fd_sc_hd__inv_2 _3181_ (.A(_2750_),
    .Y(_2751_));
 sky130_fd_sc_hd__o211ai_1 _3182_ (.A1(_2742_),
    .A2(_2748_),
    .B1(_2749_),
    .C1(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__inv_2 _3183_ (.A(\egd_top.BitStream_buffer.pc_previous[6] ),
    .Y(_2753_));
 sky130_fd_sc_hd__nand2_1 _3184_ (.A(\egd_top.BitStream_buffer.pc_previous[1] ),
    .B(\egd_top.BitStream_buffer.pc_previous[0] ),
    .Y(_2754_));
 sky130_fd_sc_hd__nand2_1 _3185_ (.A(\egd_top.BitStream_buffer.pc_previous[3] ),
    .B(\egd_top.BitStream_buffer.pc_previous[2] ),
    .Y(_2755_));
 sky130_fd_sc_hd__nand2_1 _3186_ (.A(\egd_top.BitStream_buffer.pc_previous[5] ),
    .B(\egd_top.BitStream_buffer.pc_previous[4] ),
    .Y(_2756_));
 sky130_fd_sc_hd__or3_1 _3187_ (.A(_2754_),
    .B(_2755_),
    .C(_2756_),
    .X(_2757_));
 sky130_fd_sc_hd__inv_2 _3188_ (.A(net17),
    .Y(_2758_));
 sky130_fd_sc_hd__inv_2 _3189_ (.A(net18),
    .Y(_2759_));
 sky130_fd_sc_hd__nand2_2 _3190_ (.A(_2758_),
    .B(_2759_),
    .Y(_2760_));
 sky130_fd_sc_hd__or2_1 _3191_ (.A(\egd_top.BitStream_buffer.pc_reg[0] ),
    .B(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__nand2_4 _3192_ (.A(_2760_),
    .B(\egd_top.BitStream_buffer.pc_reg[0] ),
    .Y(_2762_));
 sky130_fd_sc_hd__nand2_4 _3193_ (.A(_2761_),
    .B(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__clkinv_4 _3194_ (.A(_2763_),
    .Y(\egd_top.BitStream_buffer.pc[0] ));
 sky130_fd_sc_hd__nand2_2 _3195_ (.A(\egd_top.BitStream_buffer.pc[0] ),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2764_));
 sky130_fd_sc_hd__inv_2 _3196_ (.A(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__and3_1 _3197_ (.A(_2765_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_2766_));
 sky130_fd_sc_hd__buf_6 _3198_ (.A(_2766_),
    .X(_2767_));
 sky130_fd_sc_hd__inv_2 _3199_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2768_));
 sky130_fd_sc_hd__and3_2 _3200_ (.A(_2768_),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_2769_));
 sky130_fd_sc_hd__and2_1 _3201_ (.A(_2767_),
    .B(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__buf_6 _3202_ (.A(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__a211o_1 _3203_ (.A1(_2753_),
    .A2(_2757_),
    .B1(\egd_top.BitStream_buffer.pc[6] ),
    .C1(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__inv_2 _3204_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .Y(_2773_));
 sky130_fd_sc_hd__inv_2 _3205_ (.A(\egd_top.BitStream_buffer.buffer_index[5] ),
    .Y(_2774_));
 sky130_fd_sc_hd__inv_2 _3206_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_2775_));
 sky130_fd_sc_hd__and3_1 _3207_ (.A(_2773_),
    .B(_2774_),
    .C(_2775_),
    .X(_2776_));
 sky130_fd_sc_hd__o21ai_1 _3208_ (.A1(_2753_),
    .A2(_2776_),
    .B1(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2777_));
 sky130_fd_sc_hd__a21o_1 _3209_ (.A1(_2772_),
    .A2(_2777_),
    .B1(_2751_),
    .X(_2778_));
 sky130_fd_sc_hd__and3_1 _3210_ (.A(_2774_),
    .B(_2775_),
    .C(\egd_top.BitStream_buffer.buffer_index[6] ),
    .X(_2779_));
 sky130_fd_sc_hd__or4b_1 _3211_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(_2751_),
    .C(_2771_),
    .D_N(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__o2111ai_1 _3212_ (.A1(_2742_),
    .A2(_2748_),
    .B1(_2752_),
    .C1(_2778_),
    .D1(_2780_),
    .Y(_2781_));
 sky130_fd_sc_hd__and4_1 _3213_ (.A(_2732_),
    .B(_2739_),
    .C(net34),
    .D(net32),
    .X(_2782_));
 sky130_fd_sc_hd__nand2_1 _3214_ (.A(_2781_),
    .B(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(_2747_),
    .A1(net30),
    .S(_2783_),
    .X(_2784_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_2784_),
    .X(_0324_));
 sky130_fd_sc_hd__a21oi_1 _3217_ (.A1(_2748_),
    .A2(_2746_),
    .B1(net30),
    .Y(_2785_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(_2785_),
    .A1(net29),
    .S(_2783_),
    .X(_2786_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_2786_),
    .X(_0323_));
 sky130_fd_sc_hd__o211ai_1 _3220_ (.A1(net28),
    .A2(_2752_),
    .B1(_2778_),
    .C1(_2780_),
    .Y(_2787_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(_2787_),
    .A1(net28),
    .S(_2783_),
    .X(_2788_));
 sky130_fd_sc_hd__clkbuf_1 _3222_ (.A(_2788_),
    .X(_0322_));
 sky130_fd_sc_hd__inv_2 _3223_ (.A(net221),
    .Y(_2789_));
 sky130_fd_sc_hd__clkbuf_4 _3224_ (.A(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__nor2_1 _3225_ (.A(_2790_),
    .B(_2782_),
    .Y(_0321_));
 sky130_fd_sc_hd__buf_4 _3226_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .X(_2791_));
 sky130_fd_sc_hd__nand2_1 _3227_ (.A(_2735_),
    .B(_2734_),
    .Y(_2792_));
 sky130_fd_sc_hd__a22o_2 _3228_ (.A1(_2745_),
    .A2(_2749_),
    .B1(_2737_),
    .B2(net223),
    .X(_2793_));
 sky130_fd_sc_hd__nand2_1 _3229_ (.A(net224),
    .B(\egd_top.BitStream_buffer.buffer_index[4] ),
    .Y(_2794_));
 sky130_fd_sc_hd__or2_1 _3230_ (.A(_2774_),
    .B(_2794_),
    .X(_2795_));
 sky130_fd_sc_hd__or2_1 _3231_ (.A(_2773_),
    .B(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__buf_2 _3232_ (.A(_2796_),
    .X(_2797_));
 sky130_fd_sc_hd__buf_4 _3233_ (.A(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(net7),
    .A1(_2791_),
    .S(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__clkbuf_1 _3235_ (.A(_2799_),
    .X(_0320_));
 sky130_fd_sc_hd__buf_4 _3236_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .X(_2800_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(net6),
    .A1(_2800_),
    .S(_2798_),
    .X(_2801_));
 sky130_fd_sc_hd__clkbuf_1 _3238_ (.A(_2801_),
    .X(_0319_));
 sky130_fd_sc_hd__buf_4 _3239_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .X(_2802_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(net5),
    .A1(_2802_),
    .S(_2798_),
    .X(_2803_));
 sky130_fd_sc_hd__clkbuf_1 _3241_ (.A(_2803_),
    .X(_0318_));
 sky130_fd_sc_hd__buf_4 _3242_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .X(_2804_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(net4),
    .A1(_2804_),
    .S(_2798_),
    .X(_2805_));
 sky130_fd_sc_hd__clkbuf_1 _3244_ (.A(_2805_),
    .X(_0317_));
 sky130_fd_sc_hd__buf_4 _3245_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .X(_2806_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(net3),
    .A1(_2806_),
    .S(_2798_),
    .X(_2807_));
 sky130_fd_sc_hd__clkbuf_1 _3247_ (.A(_2807_),
    .X(_0316_));
 sky130_fd_sc_hd__buf_4 _3248_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .X(_2808_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(net2),
    .A1(_2808_),
    .S(_2798_),
    .X(_2809_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_2809_),
    .X(_0315_));
 sky130_fd_sc_hd__buf_4 _3251_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .X(_2810_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(net16),
    .A1(_2810_),
    .S(_2798_),
    .X(_2811_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_2811_),
    .X(_0314_));
 sky130_fd_sc_hd__buf_4 _3254_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .X(_2812_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(net15),
    .A1(_2812_),
    .S(_2798_),
    .X(_2813_));
 sky130_fd_sc_hd__clkbuf_1 _3256_ (.A(_2813_),
    .X(_0313_));
 sky130_fd_sc_hd__buf_4 _3257_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .X(_2814_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(net14),
    .A1(_2814_),
    .S(_2798_),
    .X(_2815_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_2815_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_8 _3260_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .X(_2816_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(net13),
    .A1(_2816_),
    .S(_2798_),
    .X(_2817_));
 sky130_fd_sc_hd__clkbuf_1 _3262_ (.A(_2817_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_8 _3263_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .X(_2818_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(net12),
    .A1(_2818_),
    .S(_2798_),
    .X(_2819_));
 sky130_fd_sc_hd__clkbuf_1 _3265_ (.A(_2819_),
    .X(_0310_));
 sky130_fd_sc_hd__buf_6 _3266_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .X(_2820_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(net11),
    .A1(_2820_),
    .S(_2797_),
    .X(_2821_));
 sky130_fd_sc_hd__clkbuf_1 _3268_ (.A(_2821_),
    .X(_0309_));
 sky130_fd_sc_hd__buf_4 _3269_ (.A(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_2822_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(net10),
    .A1(_2822_),
    .S(_2797_),
    .X(_2823_));
 sky130_fd_sc_hd__clkbuf_1 _3271_ (.A(_2823_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_8 _3272_ (.A(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_2824_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(net9),
    .A1(_2824_),
    .S(_2797_),
    .X(_2825_));
 sky130_fd_sc_hd__clkbuf_1 _3274_ (.A(_2825_),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_8 _3275_ (.A(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_2826_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(net8),
    .A1(_2826_),
    .S(_2797_),
    .X(_2827_));
 sky130_fd_sc_hd__clkbuf_1 _3277_ (.A(_2827_),
    .X(_0306_));
 sky130_fd_sc_hd__buf_4 _3278_ (.A(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_2828_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(net1),
    .A1(_2828_),
    .S(_2797_),
    .X(_2829_));
 sky130_fd_sc_hd__clkbuf_1 _3280_ (.A(_2829_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_4 _3281_ (.A(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_2830_));
 sky130_fd_sc_hd__inv_2 _3282_ (.A(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_4 _3283_ (.A(_2831_),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2832_));
 sky130_fd_sc_hd__nor2_4 _3284_ (.A(_2832_),
    .B(_2764_),
    .Y(_2833_));
 sky130_fd_sc_hd__inv_2 _3285_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_2834_));
 sky130_fd_sc_hd__inv_2 _3286_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_2835_));
 sky130_fd_sc_hd__and3_2 _3287_ (.A(_2834_),
    .B(_2835_),
    .C(\egd_top.BitStream_buffer.pc[6] ),
    .X(_2836_));
 sky130_fd_sc_hd__buf_2 _3288_ (.A(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__and2_1 _3289_ (.A(_2833_),
    .B(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3290_ (.A(_2838_),
    .X(_2839_));
 sky130_fd_sc_hd__buf_4 _3291_ (.A(_2839_),
    .X(_2840_));
 sky130_fd_sc_hd__inv_2 _3292_ (.A(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2841_));
 sky130_fd_sc_hd__nand2_4 _3293_ (.A(\egd_top.BitStream_buffer.pc[0] ),
    .B(_2841_),
    .Y(_2842_));
 sky130_fd_sc_hd__inv_2 _3294_ (.A(_2842_),
    .Y(_2843_));
 sky130_fd_sc_hd__and3_1 _3295_ (.A(_2843_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_2844_));
 sky130_fd_sc_hd__buf_4 _3296_ (.A(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__and2_1 _3297_ (.A(_2845_),
    .B(_2837_),
    .X(_2846_));
 sky130_fd_sc_hd__buf_4 _3298_ (.A(_2846_),
    .X(_2847_));
 sky130_fd_sc_hd__clkbuf_8 _3299_ (.A(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_2848_));
 sky130_fd_sc_hd__inv_2 _3300_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .Y(_2849_));
 sky130_fd_sc_hd__or3_1 _3301_ (.A(\egd_top.BitStream_buffer.pc[5] ),
    .B(_2768_),
    .C(_2834_),
    .X(_2850_));
 sky130_fd_sc_hd__inv_2 _3302_ (.A(_2850_),
    .Y(_2851_));
 sky130_fd_sc_hd__clkbuf_4 _3303_ (.A(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__nand2_1 _3304_ (.A(_2767_),
    .B(_2852_),
    .Y(_2853_));
 sky130_fd_sc_hd__clkbuf_4 _3305_ (.A(_2853_),
    .X(_2854_));
 sky130_fd_sc_hd__nand2_2 _3306_ (.A(_2763_),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2855_));
 sky130_fd_sc_hd__nor2_4 _3307_ (.A(_2832_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__and2_1 _3308_ (.A(_2856_),
    .B(_2837_),
    .X(_2857_));
 sky130_fd_sc_hd__clkbuf_4 _3309_ (.A(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__buf_4 _3310_ (.A(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_2859_));
 sky130_fd_sc_hd__nand2_1 _3311_ (.A(_2858_),
    .B(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__o21ai_1 _3312_ (.A1(_2849_),
    .A2(_2854_),
    .B1(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__a221oi_2 _3313_ (.A1(_2830_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_2848_),
    .C1(_2861_),
    .Y(_2862_));
 sky130_fd_sc_hd__buf_4 _3314_ (.A(\egd_top.BitStream_buffer.BS_buffer[25] ),
    .X(_2863_));
 sky130_fd_sc_hd__nor2_4 _3315_ (.A(_2832_),
    .B(_2842_),
    .Y(_2864_));
 sky130_fd_sc_hd__and3_2 _3316_ (.A(_2768_),
    .B(_2835_),
    .C(\egd_top.BitStream_buffer.pc[4] ),
    .X(_2865_));
 sky130_fd_sc_hd__and2_1 _3317_ (.A(_2864_),
    .B(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__clkbuf_4 _3318_ (.A(_2866_),
    .X(_2867_));
 sky130_fd_sc_hd__inv_2 _3319_ (.A(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2868_));
 sky130_fd_sc_hd__and3_1 _3320_ (.A(_2843_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__clkbuf_4 _3321_ (.A(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__and3_2 _3322_ (.A(_2768_),
    .B(_2834_),
    .C(_2835_),
    .X(_2871_));
 sky130_fd_sc_hd__clkbuf_4 _3323_ (.A(_2871_),
    .X(_2872_));
 sky130_fd_sc_hd__and2_1 _3324_ (.A(_2870_),
    .B(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__clkbuf_8 _3325_ (.A(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .X(_2874_));
 sky130_fd_sc_hd__nand2_4 _3326_ (.A(_2763_),
    .B(_2841_),
    .Y(_2875_));
 sky130_fd_sc_hd__inv_2 _3327_ (.A(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__and3_1 _3328_ (.A(_2876_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_2877_));
 sky130_fd_sc_hd__buf_4 _3329_ (.A(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__and2_1 _3330_ (.A(_2878_),
    .B(_2871_),
    .X(_2879_));
 sky130_fd_sc_hd__buf_1 _3331_ (.A(_2879_),
    .X(_2880_));
 sky130_fd_sc_hd__clkbuf_8 _3332_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .X(_2881_));
 sky130_fd_sc_hd__nand2_1 _3333_ (.A(_2880_),
    .B(_2881_),
    .Y(_2882_));
 sky130_fd_sc_hd__nand2_8 _3334_ (.A(_2831_),
    .B(_2868_),
    .Y(_2883_));
 sky130_fd_sc_hd__nor2_8 _3335_ (.A(_2883_),
    .B(_2875_),
    .Y(_2884_));
 sky130_fd_sc_hd__and2_1 _3336_ (.A(_2884_),
    .B(_2865_),
    .X(_2885_));
 sky130_fd_sc_hd__buf_1 _3337_ (.A(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__buf_4 _3338_ (.A(\egd_top.BitStream_buffer.BS_buffer[16] ),
    .X(_2887_));
 sky130_fd_sc_hd__nand2_1 _3339_ (.A(_2886_),
    .B(_2887_),
    .Y(_2888_));
 sky130_fd_sc_hd__nand2_1 _3340_ (.A(_2882_),
    .B(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__a221oi_1 _3341_ (.A1(_2863_),
    .A2(_2867_),
    .B1(_2873_),
    .B2(_2874_),
    .C1(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__inv_2 _3342_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_2891_));
 sky130_fd_sc_hd__and3_1 _3343_ (.A(_2765_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_2868_),
    .X(_2892_));
 sky130_fd_sc_hd__buf_4 _3344_ (.A(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__nand2_1 _3345_ (.A(_2893_),
    .B(_2872_),
    .Y(_2894_));
 sky130_fd_sc_hd__nor2_4 _3346_ (.A(_2883_),
    .B(_2764_),
    .Y(_2895_));
 sky130_fd_sc_hd__and2_1 _3347_ (.A(_2895_),
    .B(_2872_),
    .X(_2896_));
 sky130_fd_sc_hd__nand2_1 _3348_ (.A(_2896_),
    .B(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .Y(_2897_));
 sky130_fd_sc_hd__inv_2 _3349_ (.A(_2855_),
    .Y(_2898_));
 sky130_fd_sc_hd__and3_4 _3350_ (.A(_2898_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_2868_),
    .X(_2899_));
 sky130_fd_sc_hd__and2_1 _3351_ (.A(_2899_),
    .B(_2872_),
    .X(_2900_));
 sky130_fd_sc_hd__nand2_1 _3352_ (.A(_2900_),
    .B(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .Y(_2901_));
 sky130_fd_sc_hd__and3_4 _3353_ (.A(_2898_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(\egd_top.BitStream_buffer.pc[3] ),
    .X(_2902_));
 sky130_fd_sc_hd__and2_1 _3354_ (.A(_2902_),
    .B(_2852_),
    .X(_2903_));
 sky130_fd_sc_hd__buf_8 _3355_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .X(_2904_));
 sky130_fd_sc_hd__nand2_1 _3356_ (.A(_2903_),
    .B(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__o2111a_1 _3357_ (.A1(_2891_),
    .A2(_2894_),
    .B1(_2897_),
    .C1(_2901_),
    .D1(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__buf_4 _3358_ (.A(\egd_top.BitStream_buffer.BS_buffer[32] ),
    .X(_2907_));
 sky130_fd_sc_hd__inv_2 _3359_ (.A(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__and3_2 _3360_ (.A(_2768_),
    .B(_2834_),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_2909_));
 sky130_fd_sc_hd__clkbuf_4 _3361_ (.A(_2909_),
    .X(_2910_));
 sky130_fd_sc_hd__nand2_1 _3362_ (.A(_2884_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__clkbuf_4 _3363_ (.A(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__clkbuf_8 _3364_ (.A(\egd_top.BitStream_buffer.BS_buffer[28] ),
    .X(_2913_));
 sky130_fd_sc_hd__inv_2 _3365_ (.A(_2913_),
    .Y(_2914_));
 sky130_fd_sc_hd__clkbuf_4 _3366_ (.A(_2865_),
    .X(_2915_));
 sky130_fd_sc_hd__nand2_1 _3367_ (.A(_2878_),
    .B(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__clkbuf_4 _3368_ (.A(_2916_),
    .X(_2917_));
 sky130_fd_sc_hd__o22ai_1 _3369_ (.A1(_2908_),
    .A2(_2912_),
    .B1(_2914_),
    .B2(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__and2_1 _3370_ (.A(_2856_),
    .B(_2915_),
    .X(_2919_));
 sky130_fd_sc_hd__buf_4 _3371_ (.A(\egd_top.BitStream_buffer.BS_buffer[26] ),
    .X(_2920_));
 sky130_fd_sc_hd__and2_1 _3372_ (.A(_2833_),
    .B(_2915_),
    .X(_2921_));
 sky130_fd_sc_hd__buf_4 _3373_ (.A(\egd_top.BitStream_buffer.BS_buffer[27] ),
    .X(_2922_));
 sky130_fd_sc_hd__a22o_1 _3374_ (.A1(_2919_),
    .A2(_2920_),
    .B1(_2921_),
    .B2(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__nor2_1 _3375_ (.A(_2918_),
    .B(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__and4_1 _3376_ (.A(_2862_),
    .B(_2890_),
    .C(_2906_),
    .D(_2924_),
    .X(_2925_));
 sky130_fd_sc_hd__buf_4 _3377_ (.A(\egd_top.BitStream_buffer.BS_buffer[49] ),
    .X(_2926_));
 sky130_fd_sc_hd__nor2_8 _3378_ (.A(_2883_),
    .B(_2842_),
    .Y(_2927_));
 sky130_fd_sc_hd__and2_1 _3379_ (.A(_2927_),
    .B(_2769_),
    .X(_2928_));
 sky130_fd_sc_hd__clkbuf_2 _3380_ (.A(_2928_),
    .X(_2929_));
 sky130_fd_sc_hd__and2_2 _3381_ (.A(_2767_),
    .B(_2910_),
    .X(_2930_));
 sky130_fd_sc_hd__buf_4 _3382_ (.A(\egd_top.BitStream_buffer.BS_buffer[47] ),
    .X(_2931_));
 sky130_fd_sc_hd__and3_1 _3383_ (.A(_2876_),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .C(_2868_),
    .X(_2932_));
 sky130_fd_sc_hd__clkbuf_4 _3384_ (.A(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__and2_1 _3385_ (.A(_2933_),
    .B(_2910_),
    .X(_2934_));
 sky130_fd_sc_hd__buf_6 _3386_ (.A(\egd_top.BitStream_buffer.BS_buffer[36] ),
    .X(_2935_));
 sky130_fd_sc_hd__nand2_1 _3387_ (.A(_2934_),
    .B(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__clkbuf_4 _3388_ (.A(_2769_),
    .X(_2937_));
 sky130_fd_sc_hd__and2_1 _3389_ (.A(_2884_),
    .B(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__buf_4 _3390_ (.A(\egd_top.BitStream_buffer.BS_buffer[48] ),
    .X(_2939_));
 sky130_fd_sc_hd__nand2_1 _3391_ (.A(_2938_),
    .B(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__nand2_1 _3392_ (.A(_2936_),
    .B(_2940_),
    .Y(_2941_));
 sky130_fd_sc_hd__a221oi_2 _3393_ (.A1(_2926_),
    .A2(_2929_),
    .B1(_2930_),
    .B2(_2931_),
    .C1(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__clkbuf_8 _3394_ (.A(\egd_top.BitStream_buffer.BS_buffer[13] ),
    .X(_2943_));
 sky130_fd_sc_hd__inv_2 _3395_ (.A(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__nand2_1 _3396_ (.A(_2845_),
    .B(_2872_),
    .Y(_2945_));
 sky130_fd_sc_hd__nor2_4 _3397_ (.A(_2883_),
    .B(_2855_),
    .Y(_2946_));
 sky130_fd_sc_hd__and2_1 _3398_ (.A(_2946_),
    .B(_2872_),
    .X(_2947_));
 sky130_fd_sc_hd__nand2_1 _3399_ (.A(_2947_),
    .B(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .Y(_2948_));
 sky130_fd_sc_hd__and2_1 _3400_ (.A(_2927_),
    .B(_2872_),
    .X(_2949_));
 sky130_fd_sc_hd__nand2_1 _3401_ (.A(_2949_),
    .B(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_2950_));
 sky130_fd_sc_hd__buf_4 _3402_ (.A(\egd_top.BitStream_buffer.BS_buffer[61] ),
    .X(_2951_));
 sky130_fd_sc_hd__inv_2 _3403_ (.A(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__nand2_1 _3404_ (.A(_2845_),
    .B(_2769_),
    .Y(_2953_));
 sky130_fd_sc_hd__or2_1 _3405_ (.A(_2952_),
    .B(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__o2111a_1 _3406_ (.A1(_2944_),
    .A2(_2945_),
    .B1(_2948_),
    .C1(_2950_),
    .D1(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__and2_1 _3407_ (.A(_2933_),
    .B(_2837_),
    .X(_2956_));
 sky130_fd_sc_hd__clkbuf_8 _3408_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .X(_2957_));
 sky130_fd_sc_hd__and2_1 _3409_ (.A(_2767_),
    .B(_2837_),
    .X(_2958_));
 sky130_fd_sc_hd__clkbuf_8 _3410_ (.A(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_2959_));
 sky130_fd_sc_hd__and3_1 _3411_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .X(_2960_));
 sky130_fd_sc_hd__buf_2 _3412_ (.A(_2960_),
    .X(_2961_));
 sky130_fd_sc_hd__and2_1 _3413_ (.A(_2864_),
    .B(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__nand2_1 _3414_ (.A(_2962_),
    .B(_2816_),
    .Y(_2963_));
 sky130_fd_sc_hd__nor2_4 _3415_ (.A(_2832_),
    .B(_2875_),
    .Y(_2964_));
 sky130_fd_sc_hd__and2_1 _3416_ (.A(_2964_),
    .B(_2837_),
    .X(_2965_));
 sky130_fd_sc_hd__nand2_1 _3417_ (.A(_2965_),
    .B(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_2966_));
 sky130_fd_sc_hd__nand2_1 _3418_ (.A(_2963_),
    .B(_2966_),
    .Y(_2967_));
 sky130_fd_sc_hd__a221oi_1 _3419_ (.A1(_2956_),
    .A2(_2957_),
    .B1(_2958_),
    .B2(_2959_),
    .C1(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__and2_1 _3420_ (.A(_2933_),
    .B(_2852_),
    .X(_2969_));
 sky130_fd_sc_hd__nand2_1 _3421_ (.A(_2969_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_2970_));
 sky130_fd_sc_hd__and2_1 _3422_ (.A(_2902_),
    .B(_2837_),
    .X(_2971_));
 sky130_fd_sc_hd__nand2_1 _3423_ (.A(_2971_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_2972_));
 sky130_fd_sc_hd__and2_1 _3424_ (.A(_2964_),
    .B(_2909_),
    .X(_2973_));
 sky130_fd_sc_hd__clkbuf_8 _3425_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .X(_2974_));
 sky130_fd_sc_hd__nand2_1 _3426_ (.A(_2973_),
    .B(_2974_),
    .Y(_2975_));
 sky130_fd_sc_hd__and2_1 _3427_ (.A(_2964_),
    .B(_2852_),
    .X(_2976_));
 sky130_fd_sc_hd__nand2_1 _3428_ (.A(_2976_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_2977_));
 sky130_fd_sc_hd__and4_1 _3429_ (.A(_2970_),
    .B(_2972_),
    .C(_2975_),
    .D(_2977_),
    .X(_2978_));
 sky130_fd_sc_hd__and4_1 _3430_ (.A(_2942_),
    .B(_2955_),
    .C(_2968_),
    .D(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__clkbuf_8 _3431_ (.A(\egd_top.BitStream_buffer.BS_buffer[29] ),
    .X(_2980_));
 sky130_fd_sc_hd__inv_2 _3432_ (.A(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__nand2_1 _3433_ (.A(_2845_),
    .B(_2915_),
    .Y(_2982_));
 sky130_fd_sc_hd__or3_1 _3434_ (.A(\egd_top.BitStream_buffer.pc[4] ),
    .B(_2768_),
    .C(_2835_),
    .X(_2983_));
 sky130_fd_sc_hd__inv_2 _3435_ (.A(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__buf_2 _3436_ (.A(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__and2_1 _3437_ (.A(_2895_),
    .B(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__clkbuf_8 _3438_ (.A(\egd_top.BitStream_buffer.BS_buffer[99] ),
    .X(_2987_));
 sky130_fd_sc_hd__nand2_1 _3439_ (.A(_2986_),
    .B(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__and2_1 _3440_ (.A(_2856_),
    .B(_2985_),
    .X(_2989_));
 sky130_fd_sc_hd__clkbuf_8 _3441_ (.A(\egd_top.BitStream_buffer.BS_buffer[106] ),
    .X(_2990_));
 sky130_fd_sc_hd__nand2_1 _3442_ (.A(_2989_),
    .B(_2990_),
    .Y(_2991_));
 sky130_fd_sc_hd__and2_1 _3443_ (.A(_2946_),
    .B(_2915_),
    .X(_2992_));
 sky130_fd_sc_hd__buf_4 _3444_ (.A(\egd_top.BitStream_buffer.BS_buffer[18] ),
    .X(_2993_));
 sky130_fd_sc_hd__nand2_1 _3445_ (.A(_2992_),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__o2111a_1 _3446_ (.A1(_2981_),
    .A2(_2982_),
    .B1(_2988_),
    .C1(_2991_),
    .D1(_2994_),
    .X(_2995_));
 sky130_fd_sc_hd__buf_4 _3447_ (.A(_2961_),
    .X(_2996_));
 sky130_fd_sc_hd__and2_1 _3448_ (.A(_2893_),
    .B(_2996_),
    .X(_2997_));
 sky130_fd_sc_hd__nand2_1 _3449_ (.A(_2997_),
    .B(_2812_),
    .Y(_2998_));
 sky130_fd_sc_hd__and2_1 _3450_ (.A(_2899_),
    .B(_2996_),
    .X(_2999_));
 sky130_fd_sc_hd__nand2_1 _3451_ (.A(_2999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_3000_));
 sky130_fd_sc_hd__and2_1 _3452_ (.A(_2899_),
    .B(_2985_),
    .X(_3001_));
 sky130_fd_sc_hd__buf_4 _3453_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .X(_3002_));
 sky130_fd_sc_hd__nand2_1 _3454_ (.A(_3001_),
    .B(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__and2_1 _3455_ (.A(_2895_),
    .B(_2961_),
    .X(_3004_));
 sky130_fd_sc_hd__nand2_1 _3456_ (.A(_3004_),
    .B(_2804_),
    .Y(_3005_));
 sky130_fd_sc_hd__and4_1 _3457_ (.A(_2998_),
    .B(_3000_),
    .C(_3003_),
    .D(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__buf_4 _3458_ (.A(\egd_top.BitStream_buffer.BS_buffer[17] ),
    .X(_3007_));
 sky130_fd_sc_hd__inv_2 _3459_ (.A(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__nand2_1 _3460_ (.A(_2927_),
    .B(_2915_),
    .Y(_3009_));
 sky130_fd_sc_hd__buf_4 _3461_ (.A(\egd_top.BitStream_buffer.BS_buffer[19] ),
    .X(_3010_));
 sky130_fd_sc_hd__inv_2 _3462_ (.A(_3010_),
    .Y(_3011_));
 sky130_fd_sc_hd__nand2_1 _3463_ (.A(_2895_),
    .B(_2915_),
    .Y(_3012_));
 sky130_fd_sc_hd__o22ai_1 _3464_ (.A1(_3008_),
    .A2(_3009_),
    .B1(_3011_),
    .B2(_3012_),
    .Y(_3013_));
 sky130_fd_sc_hd__and2_1 _3465_ (.A(_2899_),
    .B(_2915_),
    .X(_3014_));
 sky130_fd_sc_hd__buf_4 _3466_ (.A(\egd_top.BitStream_buffer.BS_buffer[22] ),
    .X(_3015_));
 sky130_fd_sc_hd__and2_1 _3467_ (.A(_2893_),
    .B(_2915_),
    .X(_3016_));
 sky130_fd_sc_hd__buf_4 _3468_ (.A(\egd_top.BitStream_buffer.BS_buffer[23] ),
    .X(_3017_));
 sky130_fd_sc_hd__a22o_1 _3469_ (.A1(_3014_),
    .A2(_3015_),
    .B1(_3016_),
    .B2(_3017_),
    .X(_3018_));
 sky130_fd_sc_hd__nor2_1 _3470_ (.A(_3013_),
    .B(_3018_),
    .Y(_3019_));
 sky130_fd_sc_hd__and2_1 _3471_ (.A(_2870_),
    .B(_2996_),
    .X(_3020_));
 sky130_fd_sc_hd__nand2_1 _3472_ (.A(_3020_),
    .B(_2808_),
    .Y(_3021_));
 sky130_fd_sc_hd__and2_1 _3473_ (.A(_2927_),
    .B(_2852_),
    .X(_3022_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(_3022_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_3023_));
 sky130_fd_sc_hd__and2_1 _3475_ (.A(_2946_),
    .B(_2961_),
    .X(_3024_));
 sky130_fd_sc_hd__nand2_1 _3476_ (.A(_3024_),
    .B(_2802_),
    .Y(_3025_));
 sky130_fd_sc_hd__and2_1 _3477_ (.A(_2856_),
    .B(_2961_),
    .X(_3026_));
 sky130_fd_sc_hd__nand2_1 _3478_ (.A(_3026_),
    .B(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_3027_));
 sky130_fd_sc_hd__and4_1 _3479_ (.A(_3021_),
    .B(_3023_),
    .C(_3025_),
    .D(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__and4_1 _3480_ (.A(_2995_),
    .B(_3006_),
    .C(_3019_),
    .D(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__clkbuf_8 _3481_ (.A(\egd_top.BitStream_buffer.BS_buffer[103] ),
    .X(_3030_));
 sky130_fd_sc_hd__clkinv_4 _3482_ (.A(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__nand2_1 _3483_ (.A(_2893_),
    .B(_2985_),
    .Y(_3032_));
 sky130_fd_sc_hd__and2_1 _3484_ (.A(_2933_),
    .B(_2985_),
    .X(_3033_));
 sky130_fd_sc_hd__buf_4 _3485_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .X(_3034_));
 sky130_fd_sc_hd__nand2_1 _3486_ (.A(_3033_),
    .B(_3034_),
    .Y(_3035_));
 sky130_fd_sc_hd__and2_1 _3487_ (.A(_2964_),
    .B(_2985_),
    .X(_3036_));
 sky130_fd_sc_hd__clkbuf_8 _3488_ (.A(\egd_top.BitStream_buffer.BS_buffer[104] ),
    .X(_3037_));
 sky130_fd_sc_hd__nand2_1 _3489_ (.A(_3036_),
    .B(_3037_),
    .Y(_3038_));
 sky130_fd_sc_hd__and2_1 _3490_ (.A(_2870_),
    .B(_2915_),
    .X(_3039_));
 sky130_fd_sc_hd__buf_4 _3491_ (.A(\egd_top.BitStream_buffer.BS_buffer[21] ),
    .X(_3040_));
 sky130_fd_sc_hd__nand2_1 _3492_ (.A(_3039_),
    .B(_3040_),
    .Y(_3041_));
 sky130_fd_sc_hd__o2111a_1 _3493_ (.A1(_3031_),
    .A2(_3032_),
    .B1(_3035_),
    .C1(_3038_),
    .D1(_3041_),
    .X(_3042_));
 sky130_fd_sc_hd__and2_1 _3494_ (.A(_2833_),
    .B(_2961_),
    .X(_3043_));
 sky130_fd_sc_hd__and2_1 _3495_ (.A(_2878_),
    .B(_2961_),
    .X(_3044_));
 sky130_fd_sc_hd__a22o_1 _3496_ (.A1(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .A2(_3043_),
    .B1(_3044_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .X(_3045_));
 sky130_fd_sc_hd__nand2_1 _3497_ (.A(_2870_),
    .B(_2984_),
    .Y(_3046_));
 sky130_fd_sc_hd__inv_2 _3498_ (.A(_3046_),
    .Y(_3047_));
 sky130_fd_sc_hd__buf_4 _3499_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .X(_3048_));
 sky130_fd_sc_hd__nand2_1 _3500_ (.A(_2845_),
    .B(_2961_),
    .Y(_3049_));
 sky130_fd_sc_hd__inv_2 _3501_ (.A(_3049_),
    .Y(_3050_));
 sky130_fd_sc_hd__a22o_1 _3502_ (.A1(_3047_),
    .A2(_3048_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .B2(_3050_),
    .X(_3051_));
 sky130_fd_sc_hd__nor2_1 _3503_ (.A(_3045_),
    .B(_3051_),
    .Y(_3052_));
 sky130_fd_sc_hd__clkbuf_8 _3504_ (.A(\egd_top.BitStream_buffer.BS_buffer[105] ),
    .X(_3053_));
 sky130_fd_sc_hd__and2_1 _3505_ (.A(_2864_),
    .B(_2984_),
    .X(_3054_));
 sky130_fd_sc_hd__buf_1 _3506_ (.A(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__and2_1 _3507_ (.A(_2933_),
    .B(_2996_),
    .X(_3056_));
 sky130_fd_sc_hd__and2_1 _3508_ (.A(_2833_),
    .B(_2985_),
    .X(_3057_));
 sky130_fd_sc_hd__clkbuf_8 _3509_ (.A(\egd_top.BitStream_buffer.BS_buffer[107] ),
    .X(_3058_));
 sky130_fd_sc_hd__nand2_1 _3510_ (.A(_3057_),
    .B(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__and2_1 _3511_ (.A(_2964_),
    .B(_2961_),
    .X(_3060_));
 sky130_fd_sc_hd__nand2_1 _3512_ (.A(_3060_),
    .B(_2814_),
    .Y(_3061_));
 sky130_fd_sc_hd__nand2_1 _3513_ (.A(_3059_),
    .B(_3061_),
    .Y(_3062_));
 sky130_fd_sc_hd__a221oi_1 _3514_ (.A1(_3053_),
    .A2(_3055_),
    .B1(_3056_),
    .B2(_2806_),
    .C1(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__inv_2 _3515_ (.A(\egd_top.BitStream_buffer.BS_buffer[113] ),
    .Y(_3064_));
 sky130_fd_sc_hd__nand2_4 _3516_ (.A(_2927_),
    .B(_2996_),
    .Y(_3065_));
 sky130_fd_sc_hd__buf_4 _3517_ (.A(\egd_top.BitStream_buffer.BS_buffer[108] ),
    .X(_3066_));
 sky130_fd_sc_hd__inv_2 _3518_ (.A(_3066_),
    .Y(_3067_));
 sky130_fd_sc_hd__nand2_1 _3519_ (.A(_2878_),
    .B(_2985_),
    .Y(_3068_));
 sky130_fd_sc_hd__and2_1 _3520_ (.A(_2902_),
    .B(_2985_),
    .X(_3069_));
 sky130_fd_sc_hd__buf_4 _3521_ (.A(\egd_top.BitStream_buffer.BS_buffer[110] ),
    .X(_3070_));
 sky130_fd_sc_hd__nand2_1 _3522_ (.A(_3069_),
    .B(_3070_),
    .Y(_3071_));
 sky130_fd_sc_hd__o221a_1 _3523_ (.A1(_3064_),
    .A2(_3065_),
    .B1(_3067_),
    .B2(_3068_),
    .C1(_3071_),
    .X(_3072_));
 sky130_fd_sc_hd__and4_1 _3524_ (.A(_3042_),
    .B(_3052_),
    .C(_3063_),
    .D(_3072_),
    .X(_3073_));
 sky130_fd_sc_hd__and4_1 _3525_ (.A(_2925_),
    .B(_2979_),
    .C(_3029_),
    .D(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__inv_2 _3526_ (.A(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_3075_));
 sky130_fd_sc_hd__nand2_1 _3527_ (.A(_2870_),
    .B(_2937_),
    .Y(_3076_));
 sky130_fd_sc_hd__clkbuf_4 _3528_ (.A(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__inv_2 _3529_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .Y(_3078_));
 sky130_fd_sc_hd__nand2_1 _3530_ (.A(_2833_),
    .B(_2871_),
    .Y(_3079_));
 sky130_fd_sc_hd__buf_2 _3531_ (.A(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__or2_1 _3532_ (.A(_3078_),
    .B(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__inv_2 _3533_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_3082_));
 sky130_fd_sc_hd__nand2_1 _3534_ (.A(_2864_),
    .B(_2871_),
    .Y(_3083_));
 sky130_fd_sc_hd__buf_2 _3535_ (.A(_3083_),
    .X(_3084_));
 sky130_fd_sc_hd__or2_1 _3536_ (.A(_3082_),
    .B(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__and2_1 _3537_ (.A(_2899_),
    .B(_2937_),
    .X(_3086_));
 sky130_fd_sc_hd__clkbuf_4 _3538_ (.A(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__nand2_1 _3539_ (.A(_3087_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_3088_));
 sky130_fd_sc_hd__o2111a_1 _3540_ (.A1(_3075_),
    .A2(_3077_),
    .B1(_3081_),
    .C1(_3085_),
    .D1(_3088_),
    .X(_3089_));
 sky130_fd_sc_hd__buf_4 _3541_ (.A(\egd_top.BitStream_buffer.BS_buffer[31] ),
    .X(_3090_));
 sky130_fd_sc_hd__inv_2 _3542_ (.A(_3090_),
    .Y(_3091_));
 sky130_fd_sc_hd__nand2_1 _3543_ (.A(_2767_),
    .B(_2865_),
    .Y(_3092_));
 sky130_fd_sc_hd__clkbuf_4 _3544_ (.A(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__and2_1 _3545_ (.A(_2902_),
    .B(_2865_),
    .X(_3094_));
 sky130_fd_sc_hd__clkbuf_2 _3546_ (.A(_3094_),
    .X(_3095_));
 sky130_fd_sc_hd__buf_4 _3547_ (.A(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__clkbuf_8 _3548_ (.A(\egd_top.BitStream_buffer.BS_buffer[30] ),
    .X(_3097_));
 sky130_fd_sc_hd__nand2_1 _3549_ (.A(_3096_),
    .B(_3097_),
    .Y(_3098_));
 sky130_fd_sc_hd__and2_1 _3550_ (.A(_2856_),
    .B(_2871_),
    .X(_3099_));
 sky130_fd_sc_hd__clkbuf_4 _3551_ (.A(_3099_),
    .X(_3100_));
 sky130_fd_sc_hd__clkbuf_8 _3552_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .X(_3101_));
 sky130_fd_sc_hd__nand2_1 _3553_ (.A(_3100_),
    .B(_3101_),
    .Y(_3102_));
 sky130_fd_sc_hd__and2_2 _3554_ (.A(_2893_),
    .B(_2837_),
    .X(_3103_));
 sky130_fd_sc_hd__buf_4 _3555_ (.A(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__clkbuf_8 _3556_ (.A(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_3105_));
 sky130_fd_sc_hd__nand2_1 _3557_ (.A(_3104_),
    .B(_3105_),
    .Y(_3106_));
 sky130_fd_sc_hd__o2111a_1 _3558_ (.A1(_3091_),
    .A2(_3093_),
    .B1(_3098_),
    .C1(_3102_),
    .D1(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__inv_2 _3559_ (.A(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_3108_));
 sky130_fd_sc_hd__nand2_1 _3560_ (.A(_2893_),
    .B(_2937_),
    .Y(_3109_));
 sky130_fd_sc_hd__clkbuf_4 _3561_ (.A(_3109_),
    .X(_3110_));
 sky130_fd_sc_hd__and2_2 _3562_ (.A(_2895_),
    .B(_2769_),
    .X(_3111_));
 sky130_fd_sc_hd__buf_4 _3563_ (.A(\egd_top.BitStream_buffer.BS_buffer[51] ),
    .X(_3112_));
 sky130_fd_sc_hd__nand2_1 _3564_ (.A(_3111_),
    .B(_3112_),
    .Y(_3113_));
 sky130_fd_sc_hd__and2_1 _3565_ (.A(_2856_),
    .B(_2937_),
    .X(_3114_));
 sky130_fd_sc_hd__buf_4 _3566_ (.A(\egd_top.BitStream_buffer.BS_buffer[58] ),
    .X(_3115_));
 sky130_fd_sc_hd__nand2_1 _3567_ (.A(_3114_),
    .B(_3115_),
    .Y(_3116_));
 sky130_fd_sc_hd__and2_1 _3568_ (.A(_2933_),
    .B(_2937_),
    .X(_3117_));
 sky130_fd_sc_hd__buf_4 _3569_ (.A(_3117_),
    .X(_3118_));
 sky130_fd_sc_hd__buf_4 _3570_ (.A(\egd_top.BitStream_buffer.BS_buffer[52] ),
    .X(_3119_));
 sky130_fd_sc_hd__nand2_1 _3571_ (.A(_3118_),
    .B(_3119_),
    .Y(_3120_));
 sky130_fd_sc_hd__o2111a_1 _3572_ (.A1(_3108_),
    .A2(_3110_),
    .B1(_3113_),
    .C1(_3116_),
    .D1(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__and2_1 _3573_ (.A(_2946_),
    .B(_2909_),
    .X(_3122_));
 sky130_fd_sc_hd__buf_4 _3574_ (.A(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__clkbuf_8 _3575_ (.A(\egd_top.BitStream_buffer.BS_buffer[34] ),
    .X(_3124_));
 sky130_fd_sc_hd__and2_1 _3576_ (.A(_2927_),
    .B(_2909_),
    .X(_3125_));
 sky130_fd_sc_hd__buf_4 _3577_ (.A(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__clkbuf_8 _3578_ (.A(\egd_top.BitStream_buffer.BS_buffer[33] ),
    .X(_3127_));
 sky130_fd_sc_hd__a22o_1 _3579_ (.A1(_3123_),
    .A2(_3124_),
    .B1(_3126_),
    .B2(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__inv_2 _3580_ (.A(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_3129_));
 sky130_fd_sc_hd__nand2_1 _3581_ (.A(_2964_),
    .B(_2937_),
    .Y(_3130_));
 sky130_fd_sc_hd__clkbuf_4 _3582_ (.A(_3130_),
    .X(_3131_));
 sky130_fd_sc_hd__buf_4 _3583_ (.A(\egd_top.BitStream_buffer.BS_buffer[45] ),
    .X(_3132_));
 sky130_fd_sc_hd__inv_2 _3584_ (.A(_3132_),
    .Y(_3133_));
 sky130_fd_sc_hd__nand2_1 _3585_ (.A(_2845_),
    .B(_2910_),
    .Y(_3134_));
 sky130_fd_sc_hd__buf_4 _3586_ (.A(_3134_),
    .X(_3135_));
 sky130_fd_sc_hd__o22ai_1 _3587_ (.A1(_3129_),
    .A2(_3131_),
    .B1(_3133_),
    .B2(_3135_),
    .Y(_3136_));
 sky130_fd_sc_hd__nor2_1 _3588_ (.A(_3128_),
    .B(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__and4_1 _3589_ (.A(_3089_),
    .B(_3107_),
    .C(_3121_),
    .D(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__buf_4 _3590_ (.A(\egd_top.BitStream_buffer.BS_buffer[64] ),
    .X(_3139_));
 sky130_fd_sc_hd__and2_1 _3591_ (.A(_2884_),
    .B(_2836_),
    .X(_3140_));
 sky130_fd_sc_hd__clkbuf_2 _3592_ (.A(_3140_),
    .X(_3141_));
 sky130_fd_sc_hd__clkbuf_8 _3593_ (.A(\egd_top.BitStream_buffer.BS_buffer[63] ),
    .X(_3142_));
 sky130_fd_sc_hd__clkbuf_8 _3594_ (.A(\egd_top.BitStream_buffer.BS_buffer[42] ),
    .X(_3143_));
 sky130_fd_sc_hd__inv_2 _3595_ (.A(_3143_),
    .Y(_3144_));
 sky130_fd_sc_hd__nand2_1 _3596_ (.A(_2856_),
    .B(_2910_),
    .Y(_3145_));
 sky130_fd_sc_hd__clkbuf_8 _3597_ (.A(\egd_top.BitStream_buffer.BS_buffer[44] ),
    .X(_3146_));
 sky130_fd_sc_hd__inv_2 _3598_ (.A(_3146_),
    .Y(_3147_));
 sky130_fd_sc_hd__nand2_1 _3599_ (.A(_2878_),
    .B(_2910_),
    .Y(_3148_));
 sky130_fd_sc_hd__o22ai_1 _3600_ (.A1(_3144_),
    .A2(_3145_),
    .B1(_3147_),
    .B2(_3148_),
    .Y(_3149_));
 sky130_fd_sc_hd__a221oi_1 _3601_ (.A1(_3139_),
    .A2(_3141_),
    .B1(_2771_),
    .B2(_3142_),
    .C1(_3149_),
    .Y(_3150_));
 sky130_fd_sc_hd__inv_2 _3602_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .Y(_3151_));
 sky130_fd_sc_hd__nand2_1 _3603_ (.A(_2927_),
    .B(_2985_),
    .Y(_3152_));
 sky130_fd_sc_hd__buf_4 _3604_ (.A(\egd_top.BitStream_buffer.BS_buffer[109] ),
    .X(_3153_));
 sky130_fd_sc_hd__inv_2 _3605_ (.A(_3153_),
    .Y(_3154_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(_2845_),
    .B(_2985_),
    .Y(_3155_));
 sky130_fd_sc_hd__o22ai_1 _3607_ (.A1(_3151_),
    .A2(_3152_),
    .B1(_3154_),
    .B2(_3155_),
    .Y(_3156_));
 sky130_fd_sc_hd__and2_1 _3608_ (.A(_2884_),
    .B(_2996_),
    .X(_3157_));
 sky130_fd_sc_hd__and2_1 _3609_ (.A(_2767_),
    .B(_2985_),
    .X(_0329_));
 sky130_fd_sc_hd__buf_4 _3610_ (.A(\egd_top.BitStream_buffer.BS_buffer[111] ),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _3611_ (.A1(_2791_),
    .A2(_3157_),
    .B1(_0329_),
    .B2(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_1 _3612_ (.A(_3156_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__clkbuf_8 _3613_ (.A(\egd_top.BitStream_buffer.BS_buffer[41] ),
    .X(_0333_));
 sky130_fd_sc_hd__inv_2 _3614_ (.A(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2_1 _3615_ (.A(_2864_),
    .B(_2910_),
    .Y(_0335_));
 sky130_fd_sc_hd__clkbuf_8 _3616_ (.A(\egd_top.BitStream_buffer.BS_buffer[43] ),
    .X(_0336_));
 sky130_fd_sc_hd__inv_2 _3617_ (.A(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _3618_ (.A(_2833_),
    .B(_2910_),
    .Y(_0338_));
 sky130_fd_sc_hd__o22ai_1 _3619_ (.A1(_0334_),
    .A2(_0335_),
    .B1(_0337_),
    .B2(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__and2_1 _3620_ (.A(_2899_),
    .B(_2910_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_8 _3621_ (.A(\egd_top.BitStream_buffer.BS_buffer[38] ),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _3622_ (.A(_2893_),
    .B(_2910_),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_8 _3623_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .X(_0343_));
 sky130_fd_sc_hd__a22o_1 _3624_ (.A1(_0340_),
    .A2(_0341_),
    .B1(_0342_),
    .B2(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2_1 _3625_ (.A(_0339_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__buf_4 _3626_ (.A(\egd_top.BitStream_buffer.BS_buffer[50] ),
    .X(_0346_));
 sky130_fd_sc_hd__inv_2 _3627_ (.A(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _3628_ (.A(_2946_),
    .B(_2937_),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _3629_ (.A(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _3630_ (.A(_2902_),
    .B(_2910_),
    .Y(_0350_));
 sky130_fd_sc_hd__o22ai_1 _3631_ (.A1(_0347_),
    .A2(_0348_),
    .B1(_0349_),
    .B2(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__and2_1 _3632_ (.A(_2902_),
    .B(_2996_),
    .X(_0352_));
 sky130_fd_sc_hd__and2_1 _3633_ (.A(_2767_),
    .B(_2996_),
    .X(_0353_));
 sky130_fd_sc_hd__a22o_1 _3634_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .B1(_0353_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .X(_0354_));
 sky130_fd_sc_hd__nor2_1 _3635_ (.A(_0351_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__and4_1 _3636_ (.A(_3150_),
    .B(_0332_),
    .C(_0345_),
    .D(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__nand2_1 _3637_ (.A(_2870_),
    .B(_2852_),
    .Y(_0357_));
 sky130_fd_sc_hd__or2b_1 _3638_ (.A(_0357_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _3639_ (.A(_2946_),
    .B(_2852_),
    .X(_0359_));
 sky130_fd_sc_hd__nand2_1 _3640_ (.A(_0359_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0360_));
 sky130_fd_sc_hd__and2_1 _3641_ (.A(_2895_),
    .B(_2852_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _3642_ (.A(_0361_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0362_));
 sky130_fd_sc_hd__and2_1 _3643_ (.A(_2864_),
    .B(_2852_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _3644_ (.A(_0363_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_0364_));
 sky130_fd_sc_hd__and4_1 _3645_ (.A(_0358_),
    .B(_0360_),
    .C(_0362_),
    .D(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_4 _3646_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _3647_ (.A(_2946_),
    .B(_2836_),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _3649_ (.A(_2870_),
    .B(_2836_),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_2 _3650_ (.A(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__clkbuf_8 _3651_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_1 _3652_ (.A1(_0366_),
    .A2(_0368_),
    .B1(_0370_),
    .B2(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__and2_1 _3653_ (.A(_2899_),
    .B(_2852_),
    .X(_0373_));
 sky130_fd_sc_hd__and2_1 _3654_ (.A(_2893_),
    .B(_2852_),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _3655_ (.A1(_0373_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .B1(_0374_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0375_));
 sky130_fd_sc_hd__nor2_1 _3656_ (.A(_0372_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__and2_1 _3657_ (.A(_2870_),
    .B(_2910_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_8 _3658_ (.A(\egd_top.BitStream_buffer.BS_buffer[37] ),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _3659_ (.A(_0377_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__and2_1 _3660_ (.A(_2864_),
    .B(_2837_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_1 _3661_ (.A(_0380_),
    .B(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_0381_));
 sky130_fd_sc_hd__and2_1 _3662_ (.A(_2864_),
    .B(_2937_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _3663_ (.A(_0382_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0383_));
 sky130_fd_sc_hd__and2_1 _3664_ (.A(_2833_),
    .B(_2937_),
    .X(_0384_));
 sky130_fd_sc_hd__buf_4 _3665_ (.A(\egd_top.BitStream_buffer.BS_buffer[59] ),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _3666_ (.A(_0384_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__and4_1 _3667_ (.A(_0379_),
    .B(_0381_),
    .C(_0383_),
    .D(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__and2_1 _3668_ (.A(_2878_),
    .B(_2937_),
    .X(_0388_));
 sky130_fd_sc_hd__buf_4 _3669_ (.A(\egd_top.BitStream_buffer.BS_buffer[60] ),
    .X(_0389_));
 sky130_fd_sc_hd__nand2_1 _3670_ (.A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__and2_1 _3671_ (.A(_2902_),
    .B(_2937_),
    .X(_0391_));
 sky130_fd_sc_hd__buf_4 _3672_ (.A(\egd_top.BitStream_buffer.BS_buffer[62] ),
    .X(_0392_));
 sky130_fd_sc_hd__nand2_1 _3673_ (.A(_0391_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__and2_1 _3674_ (.A(_2895_),
    .B(_2909_),
    .X(_0394_));
 sky130_fd_sc_hd__buf_6 _3675_ (.A(\egd_top.BitStream_buffer.BS_buffer[35] ),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _3676_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__and2_1 _3677_ (.A(_2927_),
    .B(_2837_),
    .X(_0397_));
 sky130_fd_sc_hd__buf_4 _3678_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _3679_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__and4_1 _3680_ (.A(_0390_),
    .B(_0393_),
    .C(_0396_),
    .D(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__and4_1 _3681_ (.A(_0365_),
    .B(_0376_),
    .C(_0387_),
    .D(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__buf_4 _3682_ (.A(\egd_top.BitStream_buffer.BS_buffer[24] ),
    .X(_0402_));
 sky130_fd_sc_hd__inv_2 _3683_ (.A(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _3684_ (.A(_2964_),
    .B(_2915_),
    .Y(_0404_));
 sky130_fd_sc_hd__clkbuf_4 _3685_ (.A(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__buf_4 _3686_ (.A(\egd_top.BitStream_buffer.BS_buffer[20] ),
    .X(_0406_));
 sky130_fd_sc_hd__inv_2 _3687_ (.A(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(_2933_),
    .B(_2915_),
    .Y(_0408_));
 sky130_fd_sc_hd__clkbuf_4 _3689_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__o22ai_1 _3690_ (.A1(_0403_),
    .A2(_0405_),
    .B1(_0407_),
    .B2(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__and2_1 _3691_ (.A(_2902_),
    .B(_2872_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_8 _3692_ (.A(\egd_top.BitStream_buffer.BS_buffer[14] ),
    .X(_0412_));
 sky130_fd_sc_hd__and2_1 _3693_ (.A(_2767_),
    .B(_2872_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_8 _3694_ (.A(\egd_top.BitStream_buffer.BS_buffer[15] ),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _3695_ (.A1(_0411_),
    .A2(_0412_),
    .B1(_0413_),
    .B2(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__nor2_1 _3696_ (.A(_0410_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__and2_1 _3697_ (.A(_2933_),
    .B(_2872_),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _3698_ (.A(_0417_),
    .B(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0418_));
 sky130_fd_sc_hd__and2_1 _3699_ (.A(_2878_),
    .B(_2851_),
    .X(_0419_));
 sky130_fd_sc_hd__buf_6 _3700_ (.A(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _3701_ (.A(_0419_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__and2_1 _3702_ (.A(_2964_),
    .B(_2871_),
    .X(_0422_));
 sky130_fd_sc_hd__nand2_1 _3703_ (.A(_0422_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0423_));
 sky130_fd_sc_hd__and2_1 _3704_ (.A(_2884_),
    .B(_2984_),
    .X(_0424_));
 sky130_fd_sc_hd__nand2_1 _3705_ (.A(_0424_),
    .B(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_0425_));
 sky130_fd_sc_hd__and4_1 _3706_ (.A(_0418_),
    .B(_0421_),
    .C(_0423_),
    .D(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__and2_1 _3707_ (.A(_2878_),
    .B(_2836_),
    .X(_0427_));
 sky130_fd_sc_hd__buf_4 _3708_ (.A(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__nand2_1 _3709_ (.A(_0428_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_0429_));
 sky130_fd_sc_hd__and2_1 _3710_ (.A(_2899_),
    .B(_2837_),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _3711_ (.A(_0430_),
    .B(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_0431_));
 sky130_fd_sc_hd__and2_1 _3712_ (.A(_2884_),
    .B(_2851_),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_1 _3713_ (.A(_0432_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_0433_));
 sky130_fd_sc_hd__and2_1 _3714_ (.A(_2895_),
    .B(_2837_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_4 _3715_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .X(_0435_));
 sky130_fd_sc_hd__nand2_1 _3716_ (.A(_0434_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__and4_1 _3717_ (.A(_0429_),
    .B(_0431_),
    .C(_0433_),
    .D(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__and2_1 _3718_ (.A(_2856_),
    .B(_2851_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_4 _3719_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__and2_1 _3720_ (.A(_2833_),
    .B(_2851_),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_4 _3721_ (.A(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__a22o_1 _3722_ (.A1(_0439_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .B1(_0441_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_0442_));
 sky130_fd_sc_hd__buf_4 _3723_ (.A(\egd_top.BitStream_buffer.BS_buffer[98] ),
    .X(_0443_));
 sky130_fd_sc_hd__clkinv_4 _3724_ (.A(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _3725_ (.A(_2946_),
    .B(_2984_),
    .Y(_0445_));
 sky130_fd_sc_hd__clkbuf_4 _3726_ (.A(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__inv_2 _3727_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_1 _3728_ (.A(_2845_),
    .B(_2852_),
    .Y(_0448_));
 sky130_fd_sc_hd__buf_4 _3729_ (.A(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__o22ai_1 _3730_ (.A1(_0444_),
    .A2(_0446_),
    .B1(_0447_),
    .B2(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__nor2_1 _3731_ (.A(_0442_),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__and4_1 _3732_ (.A(_0416_),
    .B(_0426_),
    .C(_0437_),
    .D(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__and4_1 _3733_ (.A(_3138_),
    .B(_0356_),
    .C(_0401_),
    .D(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__o41a_1 _3734_ (.A1(\egd_top.BitStream_buffer.pc[2] ),
    .A2(\egd_top.BitStream_buffer.pc[3] ),
    .A3(\egd_top.BitStream_buffer.pc[1] ),
    .A4(\egd_top.BitStream_buffer.pc[0] ),
    .B1(_2872_),
    .X(_0454_));
 sky130_fd_sc_hd__or4_1 _3735_ (.A(\egd_top.BitStream_buffer.pc[6] ),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .C(\egd_top.BitStream_buffer.pc[5] ),
    .D(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__buf_2 _3736_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_4 _3737_ (.A(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__buf_4 _3738_ (.A(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0458_));
 sky130_fd_sc_hd__o21ai_1 _3739_ (.A1(_0458_),
    .A2(_0456_),
    .B1(_2789_),
    .Y(_0459_));
 sky130_fd_sc_hd__a31o_1 _3740_ (.A1(_3074_),
    .A2(_0453_),
    .A3(_0457_),
    .B1(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _3741_ (.A(net221),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _3742_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _3743_ (.A(_0460_),
    .B(_0462_),
    .Y(_0304_));
 sky130_fd_sc_hd__clkbuf_8 _3744_ (.A(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_8 _3745_ (.A(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_0464_));
 sky130_fd_sc_hd__inv_2 _3746_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_1 _3747_ (.A(_2858_),
    .B(_2830_),
    .Y(_0466_));
 sky130_fd_sc_hd__o21ai_1 _3748_ (.A1(_0465_),
    .A2(_2854_),
    .B1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__a221oi_2 _3749_ (.A1(_0463_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0464_),
    .C1(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__clkbuf_8 _3750_ (.A(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .X(_0469_));
 sky130_fd_sc_hd__nand2_1 _3751_ (.A(_2880_),
    .B(_2943_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _3752_ (.A(_2886_),
    .B(_3007_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_1 _3753_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__a221oi_1 _3754_ (.A1(_2920_),
    .A2(_2867_),
    .B1(_2873_),
    .B2(_0469_),
    .C1(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _3755_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _3756_ (.A(_2896_),
    .B(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _3757_ (.A(_2900_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_0476_));
 sky130_fd_sc_hd__clkbuf_8 _3758_ (.A(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .X(_0477_));
 sky130_fd_sc_hd__nand2_1 _3759_ (.A(_2903_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__o2111a_1 _3760_ (.A1(_0474_),
    .A2(_2894_),
    .B1(_0475_),
    .C1(_0476_),
    .D1(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__inv_2 _3761_ (.A(_3127_),
    .Y(_0480_));
 sky130_fd_sc_hd__o22ai_1 _3762_ (.A1(_0480_),
    .A2(_2912_),
    .B1(_2981_),
    .B2(_2917_),
    .Y(_0481_));
 sky130_fd_sc_hd__a22o_1 _3763_ (.A1(_2919_),
    .A2(_2922_),
    .B1(_2921_),
    .B2(_2913_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_1 _3764_ (.A(_0481_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__and4_1 _3765_ (.A(_0468_),
    .B(_0473_),
    .C(_0479_),
    .D(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__nand2_1 _3766_ (.A(_2934_),
    .B(_0378_),
    .Y(_0485_));
 sky130_fd_sc_hd__nand2_1 _3767_ (.A(_2938_),
    .B(_2926_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand2_1 _3768_ (.A(_0485_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__a221oi_2 _3769_ (.A1(_0346_),
    .A2(_2929_),
    .B1(_2930_),
    .B2(_2939_),
    .C1(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _3770_ (.A(_0412_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _3771_ (.A(_2947_),
    .B(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _3772_ (.A(_2949_),
    .B(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_2 _3773_ (.A(_0392_),
    .Y(_0492_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(_0492_),
    .B(_2953_),
    .X(_0493_));
 sky130_fd_sc_hd__o2111a_1 _3775_ (.A1(_0489_),
    .A2(_2945_),
    .B1(_0490_),
    .C1(_0491_),
    .D1(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__buf_4 _3776_ (.A(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_0495_));
 sky130_fd_sc_hd__nand2_1 _3777_ (.A(_2962_),
    .B(_2818_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _3778_ (.A(_2965_),
    .B(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .Y(_0497_));
 sky130_fd_sc_hd__nand2_1 _3779_ (.A(_0496_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__a221oi_1 _3780_ (.A1(_2956_),
    .A2(_0371_),
    .B1(_2958_),
    .B2(_0495_),
    .C1(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _3781_ (.A(_2969_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _3782_ (.A(_2971_),
    .B(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .Y(_0501_));
 sky130_fd_sc_hd__nand2_1 _3783_ (.A(_2973_),
    .B(_0333_),
    .Y(_0502_));
 sky130_fd_sc_hd__nand2_1 _3784_ (.A(_2976_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_0503_));
 sky130_fd_sc_hd__and4_1 _3785_ (.A(_0500_),
    .B(_0501_),
    .C(_0502_),
    .D(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__and4_1 _3786_ (.A(_0488_),
    .B(_0494_),
    .C(_0499_),
    .D(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__inv_2 _3787_ (.A(_3097_),
    .Y(_0506_));
 sky130_fd_sc_hd__nand2_1 _3788_ (.A(_2986_),
    .B(_3034_),
    .Y(_0507_));
 sky130_fd_sc_hd__nand2_1 _3789_ (.A(_2989_),
    .B(_3058_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_1 _3790_ (.A(_2992_),
    .B(_3010_),
    .Y(_0509_));
 sky130_fd_sc_hd__o2111a_1 _3791_ (.A1(_0506_),
    .A2(_2982_),
    .B1(_0507_),
    .C1(_0508_),
    .D1(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _3792_ (.A(_2997_),
    .B(_2814_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _3793_ (.A(_2999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_0512_));
 sky130_fd_sc_hd__nand2_1 _3794_ (.A(_3001_),
    .B(_3030_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _3795_ (.A(_3004_),
    .B(_2806_),
    .Y(_0514_));
 sky130_fd_sc_hd__and4_1 _3796_ (.A(_0511_),
    .B(_0512_),
    .C(_0513_),
    .D(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__inv_2 _3797_ (.A(_2993_),
    .Y(_0516_));
 sky130_fd_sc_hd__o22ai_1 _3798_ (.A1(_0516_),
    .A2(_3009_),
    .B1(_0407_),
    .B2(_3012_),
    .Y(_0517_));
 sky130_fd_sc_hd__a22o_1 _3799_ (.A1(_3014_),
    .A2(_3017_),
    .B1(_3016_),
    .B2(_0402_),
    .X(_0518_));
 sky130_fd_sc_hd__nor2_1 _3800_ (.A(_0517_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_1 _3801_ (.A(_3020_),
    .B(_2810_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _3802_ (.A(_3022_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _3803_ (.A(_3024_),
    .B(_2804_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _3804_ (.A(_3026_),
    .B(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_0523_));
 sky130_fd_sc_hd__and4_1 _3805_ (.A(_0520_),
    .B(_0521_),
    .C(_0522_),
    .D(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__and4_1 _3806_ (.A(_0510_),
    .B(_0515_),
    .C(_0519_),
    .D(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__clkinv_4 _3807_ (.A(_3037_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_1 _3808_ (.A(_3033_),
    .B(_3048_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _3809_ (.A(_3036_),
    .B(_3053_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_1 _3810_ (.A(_3039_),
    .B(_3015_),
    .Y(_0529_));
 sky130_fd_sc_hd__o2111a_1 _3811_ (.A1(_0526_),
    .A2(_3032_),
    .B1(_0527_),
    .C1(_0528_),
    .D1(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _3812_ (.A1(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .A2(_3043_),
    .B1(_3044_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _3813_ (.A1(_3047_),
    .A2(_3002_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .B2(_3050_),
    .X(_0532_));
 sky130_fd_sc_hd__nor2_1 _3814_ (.A(_0531_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_1 _3815_ (.A(_3057_),
    .B(_3066_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _3816_ (.A(_3060_),
    .B(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_0535_));
 sky130_fd_sc_hd__nand2_1 _3817_ (.A(_0534_),
    .B(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__a221oi_1 _3818_ (.A1(_2990_),
    .A2(_3055_),
    .B1(_3056_),
    .B2(_2808_),
    .C1(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__inv_2 _3819_ (.A(\egd_top.BitStream_buffer.BS_buffer[114] ),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _3820_ (.A(_3069_),
    .B(_0330_),
    .Y(_0539_));
 sky130_fd_sc_hd__o221a_1 _3821_ (.A1(_0538_),
    .A2(_3065_),
    .B1(_3154_),
    .B2(_3068_),
    .C1(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__and4_1 _3822_ (.A(_0530_),
    .B(_0533_),
    .C(_0537_),
    .D(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__and4_1 _3823_ (.A(_0484_),
    .B(_0505_),
    .C(_0525_),
    .D(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__inv_2 _3824_ (.A(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0543_));
 sky130_fd_sc_hd__inv_2 _3825_ (.A(\egd_top.BitStream_buffer.BS_buffer[12] ),
    .Y(_0544_));
 sky130_fd_sc_hd__or2_1 _3826_ (.A(_0544_),
    .B(_3080_),
    .X(_0545_));
 sky130_fd_sc_hd__inv_2 _3827_ (.A(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0546_));
 sky130_fd_sc_hd__or2_1 _3828_ (.A(_0546_),
    .B(_3084_),
    .X(_0547_));
 sky130_fd_sc_hd__nand2_1 _3829_ (.A(_3087_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_0548_));
 sky130_fd_sc_hd__o2111a_1 _3830_ (.A1(_0543_),
    .A2(_3077_),
    .B1(_0545_),
    .C1(_0547_),
    .D1(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_1 _3831_ (.A(_3096_),
    .B(_3090_),
    .Y(_0550_));
 sky130_fd_sc_hd__clkbuf_8 _3832_ (.A(\egd_top.BitStream_buffer.BS_buffer[11] ),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _3833_ (.A(_3100_),
    .B(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__clkbuf_8 _3834_ (.A(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_1 _3835_ (.A(_3104_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__o2111a_1 _3836_ (.A1(_2908_),
    .A2(_3093_),
    .B1(_0550_),
    .C1(_0552_),
    .D1(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _3837_ (.A(_3111_),
    .B(_3119_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _3838_ (.A(_3114_),
    .B(_0385_),
    .Y(_0557_));
 sky130_fd_sc_hd__nand2_1 _3839_ (.A(_3118_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_0558_));
 sky130_fd_sc_hd__o2111a_1 _3840_ (.A1(_3129_),
    .A2(_3110_),
    .B1(_0556_),
    .C1(_0557_),
    .D1(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _3841_ (.A1(_3123_),
    .A2(_0395_),
    .B1(_3126_),
    .B2(_3124_),
    .X(_0560_));
 sky130_fd_sc_hd__inv_2 _3842_ (.A(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0561_));
 sky130_fd_sc_hd__o22ai_1 _3843_ (.A1(_0561_),
    .A2(_3131_),
    .B1(_0349_),
    .B2(_3135_),
    .Y(_0562_));
 sky130_fd_sc_hd__nor2_1 _3844_ (.A(_0560_),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__and4_1 _3845_ (.A(_0549_),
    .B(_0555_),
    .C(_0559_),
    .D(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__o22ai_1 _3846_ (.A1(_0337_),
    .A2(_3145_),
    .B1(_3133_),
    .B2(_3148_),
    .Y(_0565_));
 sky130_fd_sc_hd__a221oi_1 _3847_ (.A1(_0398_),
    .A2(_3141_),
    .B1(_2771_),
    .B2(_3139_),
    .C1(_0565_),
    .Y(_0566_));
 sky130_fd_sc_hd__inv_2 _3848_ (.A(_3070_),
    .Y(_0567_));
 sky130_fd_sc_hd__o22ai_1 _3849_ (.A1(_0444_),
    .A2(_3152_),
    .B1(_0567_),
    .B2(_3155_),
    .Y(_0568_));
 sky130_fd_sc_hd__a22o_1 _3850_ (.A1(_2800_),
    .A2(_3157_),
    .B1(_0329_),
    .B2(_2791_),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_1 _3851_ (.A(_0568_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__o22ai_1 _3852_ (.A1(_3144_),
    .A2(_0335_),
    .B1(_3147_),
    .B2(_0338_),
    .Y(_0571_));
 sky130_fd_sc_hd__a22o_1 _3853_ (.A1(_0340_),
    .A2(_0343_),
    .B1(_0342_),
    .B2(_2974_),
    .X(_0572_));
 sky130_fd_sc_hd__nor2_1 _3854_ (.A(_0571_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__inv_2 _3855_ (.A(_3112_),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_2 _3856_ (.A(_2931_),
    .Y(_0575_));
 sky130_fd_sc_hd__o22ai_1 _3857_ (.A1(_0574_),
    .A2(_0348_),
    .B1(_0575_),
    .B2(_0350_),
    .Y(_0576_));
 sky130_fd_sc_hd__a22o_1 _3858_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .B1(_0353_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .X(_0577_));
 sky130_fd_sc_hd__nor2_1 _3859_ (.A(_0576_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__and4_1 _3860_ (.A(_0566_),
    .B(_0570_),
    .C(_0573_),
    .D(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__or2b_1 _3861_ (.A(_0357_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_1 _3862_ (.A(_0359_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _3863_ (.A(_0361_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0582_));
 sky130_fd_sc_hd__clkbuf_8 _3864_ (.A(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _3865_ (.A(_0363_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__and4_1 _3866_ (.A(_0580_),
    .B(_0581_),
    .C(_0582_),
    .D(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__a22o_1 _3867_ (.A1(_0435_),
    .A2(_0368_),
    .B1(_0370_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_0586_));
 sky130_fd_sc_hd__buf_4 _3868_ (.A(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _3869_ (.A1(_0373_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .B1(_0374_),
    .B2(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__nor2_1 _3870_ (.A(_0586_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__nand2_1 _3871_ (.A(_0377_),
    .B(_0341_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _3872_ (.A(_0380_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _3873_ (.A(_0382_),
    .B(_3115_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand2_1 _3874_ (.A(_0384_),
    .B(_0389_),
    .Y(_0593_));
 sky130_fd_sc_hd__and4_1 _3875_ (.A(_0590_),
    .B(_0591_),
    .C(_0592_),
    .D(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__nand2_1 _3876_ (.A(_0388_),
    .B(_2951_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(_0391_),
    .B(_3142_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _3878_ (.A(_0394_),
    .B(_2935_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _3879_ (.A(_0397_),
    .B(_0366_),
    .Y(_0598_));
 sky130_fd_sc_hd__and4_1 _3880_ (.A(_0595_),
    .B(_0596_),
    .C(_0597_),
    .D(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__and4_2 _3881_ (.A(_0585_),
    .B(_0589_),
    .C(_0594_),
    .D(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__inv_2 _3882_ (.A(_2863_),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_2 _3883_ (.A(_3040_),
    .Y(_0602_));
 sky130_fd_sc_hd__o22ai_1 _3884_ (.A1(_0601_),
    .A2(_0405_),
    .B1(_0602_),
    .B2(_0409_),
    .Y(_0603_));
 sky130_fd_sc_hd__a22o_1 _3885_ (.A1(_0411_),
    .A2(_0414_),
    .B1(_0413_),
    .B2(_2887_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _3886_ (.A(_0603_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__nand2_1 _3887_ (.A(_0417_),
    .B(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .Y(_0606_));
 sky130_fd_sc_hd__buf_8 _3888_ (.A(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_1 _3889_ (.A(_0419_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _3890_ (.A(_0422_),
    .B(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .Y(_0609_));
 sky130_fd_sc_hd__buf_4 _3891_ (.A(\egd_top.BitStream_buffer.BS_buffer[97] ),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_1 _3892_ (.A(_0424_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__and4_1 _3893_ (.A(_0606_),
    .B(_0608_),
    .C(_0609_),
    .D(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__nand2_1 _3894_ (.A(_0428_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_0613_));
 sky130_fd_sc_hd__nand2_1 _3895_ (.A(_0430_),
    .B(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_1 _3896_ (.A(_0432_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_1 _3897_ (.A(_0434_),
    .B(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_0616_));
 sky130_fd_sc_hd__and4_1 _3898_ (.A(_0613_),
    .B(_0614_),
    .C(_0615_),
    .D(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__a22o_1 _3899_ (.A1(_0439_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .B1(_0441_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_0618_));
 sky130_fd_sc_hd__clkinv_4 _3900_ (.A(_2987_),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_2 _3901_ (.A(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_0620_));
 sky130_fd_sc_hd__o22ai_1 _3902_ (.A1(_0619_),
    .A2(_0446_),
    .B1(_0620_),
    .B2(_0449_),
    .Y(_0621_));
 sky130_fd_sc_hd__nor2_1 _3903_ (.A(_0618_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__and4_1 _3904_ (.A(_0605_),
    .B(_0612_),
    .C(_0617_),
    .D(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__and4_1 _3905_ (.A(_0564_),
    .B(_0579_),
    .C(_0600_),
    .D(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__buf_4 _3906_ (.A(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0625_));
 sky130_fd_sc_hd__o21ai_1 _3907_ (.A1(_0625_),
    .A2(_0456_),
    .B1(_2789_),
    .Y(_0626_));
 sky130_fd_sc_hd__a31o_1 _3908_ (.A1(_0542_),
    .A2(_0624_),
    .A3(_0457_),
    .B1(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__nand2_1 _3909_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_0627_),
    .B(_0628_),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_1 _3911_ (.A(_2870_),
    .B(_2872_),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _3912_ (.A(_2866_),
    .B(_2922_),
    .Y(_0630_));
 sky130_fd_sc_hd__o21ai_1 _3913_ (.A1(_2891_),
    .A2(_0629_),
    .B1(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__a221oi_1 _3914_ (.A1(_0412_),
    .A2(_2880_),
    .B1(_2993_),
    .B2(_2886_),
    .C1(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand2_1 _3915_ (.A(_2857_),
    .B(_0463_),
    .Y(_0633_));
 sky130_fd_sc_hd__o21ai_1 _3916_ (.A1(_3151_),
    .A2(_2853_),
    .B1(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__a221oi_2 _3917_ (.A1(_2848_),
    .A2(_2839_),
    .B1(_2846_),
    .B2(_2959_),
    .C1(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2_1 _3918_ (.A(_2896_),
    .B(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_1 _3919_ (.A(_2900_),
    .B(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .Y(_0637_));
 sky130_fd_sc_hd__buf_4 _3920_ (.A(\egd_top.BitStream_buffer.BS_buffer[96] ),
    .X(_0638_));
 sky130_fd_sc_hd__nand2_1 _3921_ (.A(_2903_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__o2111a_1 _3922_ (.A1(_3082_),
    .A2(_2894_),
    .B1(_0636_),
    .C1(_0637_),
    .D1(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__inv_2 _3923_ (.A(_3124_),
    .Y(_0641_));
 sky130_fd_sc_hd__o22ai_1 _3924_ (.A1(_0641_),
    .A2(_2912_),
    .B1(_0506_),
    .B2(_2917_),
    .Y(_0642_));
 sky130_fd_sc_hd__a22o_1 _3925_ (.A1(_2919_),
    .A2(_2913_),
    .B1(_2921_),
    .B2(_2980_),
    .X(_0643_));
 sky130_fd_sc_hd__nor2_1 _3926_ (.A(_0642_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__and4_1 _3927_ (.A(_0632_),
    .B(_0635_),
    .C(_0640_),
    .D(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nand2_1 _3928_ (.A(_2934_),
    .B(_0341_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _3929_ (.A(_2938_),
    .B(_0346_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _3930_ (.A(_0646_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__a221oi_2 _3931_ (.A1(_3112_),
    .A2(_2929_),
    .B1(_2930_),
    .B2(_2926_),
    .C1(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__inv_2 _3932_ (.A(_0414_),
    .Y(_0650_));
 sky130_fd_sc_hd__nand2_1 _3933_ (.A(_2947_),
    .B(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .Y(_0651_));
 sky130_fd_sc_hd__nand2_1 _3934_ (.A(_2949_),
    .B(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _3935_ (.A(_3142_),
    .Y(_0653_));
 sky130_fd_sc_hd__or2_1 _3936_ (.A(_0653_),
    .B(_2953_),
    .X(_0654_));
 sky130_fd_sc_hd__o2111a_1 _3937_ (.A1(_0650_),
    .A2(_2945_),
    .B1(_0651_),
    .C1(_0652_),
    .D1(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__clkbuf_8 _3938_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .X(_0656_));
 sky130_fd_sc_hd__buf_4 _3939_ (.A(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .X(_0657_));
 sky130_fd_sc_hd__nand2_1 _3940_ (.A(_2962_),
    .B(_2820_),
    .Y(_0658_));
 sky130_fd_sc_hd__nand2_1 _3941_ (.A(_2965_),
    .B(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .Y(_0659_));
 sky130_fd_sc_hd__nand2_1 _3942_ (.A(_0658_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__a221oi_1 _3943_ (.A1(_2956_),
    .A2(_0656_),
    .B1(_2958_),
    .B2(_0657_),
    .C1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(_2969_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_0662_));
 sky130_fd_sc_hd__nand2_1 _3945_ (.A(_2971_),
    .B(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _3946_ (.A(_2973_),
    .B(_3143_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _3947_ (.A(_2976_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_0665_));
 sky130_fd_sc_hd__and4_1 _3948_ (.A(_0662_),
    .B(_0663_),
    .C(_0664_),
    .D(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__and4_1 _3949_ (.A(_0649_),
    .B(_0655_),
    .C(_0661_),
    .D(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__nand2_1 _3950_ (.A(_2986_),
    .B(_3048_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_1 _3951_ (.A(_2989_),
    .B(_3066_),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _3952_ (.A(_2992_),
    .B(_0406_),
    .Y(_0670_));
 sky130_fd_sc_hd__o2111a_1 _3953_ (.A1(_3091_),
    .A2(_2982_),
    .B1(_0668_),
    .C1(_0669_),
    .D1(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_1 _3954_ (.A(_2997_),
    .B(_2816_),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2_1 _3955_ (.A(_2999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_0673_));
 sky130_fd_sc_hd__nand2_1 _3956_ (.A(_3001_),
    .B(_3037_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _3957_ (.A(_3004_),
    .B(_2808_),
    .Y(_0675_));
 sky130_fd_sc_hd__and4_1 _3958_ (.A(_0672_),
    .B(_0673_),
    .C(_0674_),
    .D(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__o22ai_1 _3959_ (.A1(_3011_),
    .A2(_3009_),
    .B1(_0602_),
    .B2(_3012_),
    .Y(_0677_));
 sky130_fd_sc_hd__a22o_1 _3960_ (.A1(_3014_),
    .A2(_0402_),
    .B1(_3016_),
    .B2(_2863_),
    .X(_0678_));
 sky130_fd_sc_hd__nor2_1 _3961_ (.A(_0677_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__nand2_1 _3962_ (.A(_3020_),
    .B(_2812_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _3963_ (.A(_3022_),
    .B(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _3964_ (.A(_3024_),
    .B(_2806_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _3965_ (.A(_3026_),
    .B(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_0683_));
 sky130_fd_sc_hd__and4_1 _3966_ (.A(_0680_),
    .B(_0681_),
    .C(_0682_),
    .D(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__and4_1 _3967_ (.A(_0671_),
    .B(_0676_),
    .C(_0679_),
    .D(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__clkinv_4 _3968_ (.A(_3053_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _3969_ (.A(_3033_),
    .B(_3002_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(_3036_),
    .B(_2990_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2_1 _3971_ (.A(_3039_),
    .B(_3017_),
    .Y(_0689_));
 sky130_fd_sc_hd__o2111a_1 _3972_ (.A1(_0686_),
    .A2(_3032_),
    .B1(_0687_),
    .C1(_0688_),
    .D1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__a22o_1 _3973_ (.A1(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .A2(_3043_),
    .B1(_3044_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .X(_0691_));
 sky130_fd_sc_hd__a22o_1 _3974_ (.A1(_3047_),
    .A2(_3030_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .B2(_3050_),
    .X(_0692_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_0691_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__nand2_1 _3976_ (.A(_3057_),
    .B(_3153_),
    .Y(_0694_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(_3060_),
    .B(_2818_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _3978_ (.A(_0694_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__a221oi_1 _3979_ (.A1(_3058_),
    .A2(_3055_),
    .B1(_3056_),
    .B2(_2810_),
    .C1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__inv_2 _3980_ (.A(\egd_top.BitStream_buffer.BS_buffer[115] ),
    .Y(_0698_));
 sky130_fd_sc_hd__nand2_1 _3981_ (.A(_3069_),
    .B(_2791_),
    .Y(_0699_));
 sky130_fd_sc_hd__o221a_1 _3982_ (.A1(_0698_),
    .A2(_3065_),
    .B1(_0567_),
    .B2(_3068_),
    .C1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__and4_1 _3983_ (.A(_0690_),
    .B(_0693_),
    .C(_0697_),
    .D(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__and4_1 _3984_ (.A(_0645_),
    .B(_0667_),
    .C(_0685_),
    .D(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__or2_1 _3985_ (.A(_2944_),
    .B(_3080_),
    .X(_0703_));
 sky130_fd_sc_hd__or2_1 _3986_ (.A(_3078_),
    .B(_3084_),
    .X(_0704_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(_3087_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_0705_));
 sky130_fd_sc_hd__o2111a_1 _3988_ (.A1(_3108_),
    .A2(_3077_),
    .B1(_0703_),
    .C1(_0704_),
    .D1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__nand2_1 _3989_ (.A(_3096_),
    .B(_2907_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand2_1 _3990_ (.A(_3100_),
    .B(_2881_),
    .Y(_0708_));
 sky130_fd_sc_hd__buf_4 _3991_ (.A(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_0709_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(_3104_),
    .B(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__o2111a_1 _3993_ (.A1(_0480_),
    .A2(_3093_),
    .B1(_0707_),
    .C1(_0708_),
    .D1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__nand2_1 _3994_ (.A(_3111_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_0712_));
 sky130_fd_sc_hd__nand2_1 _3995_ (.A(_3114_),
    .B(_0389_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _3996_ (.A(_3118_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_0714_));
 sky130_fd_sc_hd__o2111a_1 _3997_ (.A1(_0561_),
    .A2(_3110_),
    .B1(_0712_),
    .C1(_0713_),
    .D1(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__a22o_1 _3998_ (.A1(_3123_),
    .A2(_2935_),
    .B1(_3126_),
    .B2(_0395_),
    .X(_0716_));
 sky130_fd_sc_hd__inv_2 _3999_ (.A(_3115_),
    .Y(_0717_));
 sky130_fd_sc_hd__o22ai_1 _4000_ (.A1(_0717_),
    .A2(_3131_),
    .B1(_0575_),
    .B2(_3135_),
    .Y(_0718_));
 sky130_fd_sc_hd__nor2_1 _4001_ (.A(_0716_),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__and4_1 _4002_ (.A(_0706_),
    .B(_0711_),
    .C(_0715_),
    .D(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__o22ai_1 _4003_ (.A1(_3147_),
    .A2(_3145_),
    .B1(_0349_),
    .B2(_3148_),
    .Y(_0721_));
 sky130_fd_sc_hd__a221oi_1 _4004_ (.A1(_0366_),
    .A2(_3141_),
    .B1(_2771_),
    .B2(_0398_),
    .C1(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__inv_2 _4005_ (.A(_0330_),
    .Y(_0723_));
 sky130_fd_sc_hd__o22ai_1 _4006_ (.A1(_0619_),
    .A2(_3152_),
    .B1(_0723_),
    .B2(_3155_),
    .Y(_0724_));
 sky130_fd_sc_hd__a22o_1 _4007_ (.A1(_2802_),
    .A2(_3157_),
    .B1(_0329_),
    .B2(_2800_),
    .X(_0725_));
 sky130_fd_sc_hd__nor2_1 _4008_ (.A(_0724_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__o22ai_1 _4009_ (.A1(_0337_),
    .A2(_0335_),
    .B1(_3133_),
    .B2(_0338_),
    .Y(_0727_));
 sky130_fd_sc_hd__a22o_1 _4010_ (.A1(_0340_),
    .A2(_2974_),
    .B1(_0342_),
    .B2(_0333_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _4011_ (.A(_0727_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__inv_2 _4012_ (.A(_3119_),
    .Y(_0730_));
 sky130_fd_sc_hd__inv_2 _4013_ (.A(_2939_),
    .Y(_0731_));
 sky130_fd_sc_hd__o22ai_1 _4014_ (.A1(_0730_),
    .A2(_0348_),
    .B1(_0731_),
    .B2(_0350_),
    .Y(_0732_));
 sky130_fd_sc_hd__a22o_1 _4015_ (.A1(_0352_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .B1(_0353_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .X(_0733_));
 sky130_fd_sc_hd__nor2_1 _4016_ (.A(_0732_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__and4_1 _4017_ (.A(_0722_),
    .B(_0726_),
    .C(_0729_),
    .D(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__or2b_1 _4018_ (.A(_0357_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(_0359_),
    .B(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(_0361_),
    .B(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _4021_ (.A(_0363_),
    .B(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .Y(_0739_));
 sky130_fd_sc_hd__and4_1 _4022_ (.A(_0736_),
    .B(_0737_),
    .C(_0738_),
    .D(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _4023_ (.A1(_2957_),
    .A2(_0368_),
    .B1(_0370_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_0741_));
 sky130_fd_sc_hd__clkbuf_8 _4024_ (.A(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_0742_));
 sky130_fd_sc_hd__a22o_1 _4025_ (.A1(_0373_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .B1(_0374_),
    .B2(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__nor2_1 _4026_ (.A(_0741_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__nand2_1 _4027_ (.A(_0377_),
    .B(_0343_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand2_1 _4028_ (.A(_0380_),
    .B(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(_0382_),
    .B(_0385_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _4030_ (.A(_0384_),
    .B(_2951_),
    .Y(_0748_));
 sky130_fd_sc_hd__and4_1 _4031_ (.A(_0745_),
    .B(_0746_),
    .C(_0747_),
    .D(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__nand2_1 _4032_ (.A(_0388_),
    .B(_0392_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2_1 _4033_ (.A(_0391_),
    .B(_3139_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _4034_ (.A(_0394_),
    .B(_0378_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _4035_ (.A(_0397_),
    .B(_0435_),
    .Y(_0753_));
 sky130_fd_sc_hd__and4_1 _4036_ (.A(_0750_),
    .B(_0751_),
    .C(_0752_),
    .D(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__and4_1 _4037_ (.A(_0740_),
    .B(_0744_),
    .C(_0749_),
    .D(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__inv_2 _4038_ (.A(_2920_),
    .Y(_0756_));
 sky130_fd_sc_hd__inv_2 _4039_ (.A(_3015_),
    .Y(_0757_));
 sky130_fd_sc_hd__o22ai_1 _4040_ (.A1(_0756_),
    .A2(_0405_),
    .B1(_0757_),
    .B2(_0409_),
    .Y(_0758_));
 sky130_fd_sc_hd__a22o_1 _4041_ (.A1(_0411_),
    .A2(_2887_),
    .B1(_0413_),
    .B2(_3007_),
    .X(_0759_));
 sky130_fd_sc_hd__nor2_1 _4042_ (.A(_0758_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(_0417_),
    .B(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .Y(_0761_));
 sky130_fd_sc_hd__nand2_1 _4044_ (.A(_0419_),
    .B(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_1 _4045_ (.A(_0422_),
    .B(\egd_top.BitStream_buffer.BS_buffer[10] ),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(_0424_),
    .B(_0443_),
    .Y(_0764_));
 sky130_fd_sc_hd__and4_1 _4047_ (.A(_0761_),
    .B(_0762_),
    .C(_0763_),
    .D(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__nand2_1 _4048_ (.A(_0428_),
    .B(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .Y(_0766_));
 sky130_fd_sc_hd__nand2_1 _4049_ (.A(_0430_),
    .B(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .Y(_0767_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(_0432_),
    .B(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .Y(_0768_));
 sky130_fd_sc_hd__nand2_1 _4051_ (.A(_0434_),
    .B(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_0769_));
 sky130_fd_sc_hd__and4_1 _4052_ (.A(_0766_),
    .B(_0767_),
    .C(_0768_),
    .D(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _4053_ (.A1(_0439_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .B1(_0441_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .X(_0771_));
 sky130_fd_sc_hd__inv_2 _4054_ (.A(\egd_top.BitStream_buffer.BS_buffer[100] ),
    .Y(_0772_));
 sky130_fd_sc_hd__o22ai_1 _4055_ (.A1(_0772_),
    .A2(_0446_),
    .B1(_2849_),
    .B2(_0449_),
    .Y(_0773_));
 sky130_fd_sc_hd__nor2_1 _4056_ (.A(_0771_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__and4_1 _4057_ (.A(_0760_),
    .B(_0765_),
    .C(_0770_),
    .D(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__and4_1 _4058_ (.A(_0720_),
    .B(_0735_),
    .C(_0755_),
    .D(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__buf_4 _4059_ (.A(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .X(_0777_));
 sky130_fd_sc_hd__o21ai_1 _4060_ (.A1(_0777_),
    .A2(_0456_),
    .B1(_2789_),
    .Y(_0778_));
 sky130_fd_sc_hd__a31o_1 _4061_ (.A1(_0702_),
    .A2(_0776_),
    .A3(_0457_),
    .B1(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__nand2_1 _4062_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_0780_));
 sky130_fd_sc_hd__nand2_1 _4063_ (.A(_0779_),
    .B(_0780_),
    .Y(_0302_));
 sky130_fd_sc_hd__clkbuf_4 _4064_ (.A(_3050_),
    .X(_0781_));
 sky130_fd_sc_hd__clkbuf_4 _4065_ (.A(_3047_),
    .X(_0782_));
 sky130_fd_sc_hd__clkbuf_4 _4066_ (.A(_3043_),
    .X(_0783_));
 sky130_fd_sc_hd__clkbuf_4 _4067_ (.A(_3044_),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _4068_ (.A1(\egd_top.BitStream_buffer.BS_buffer[126] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_2828_),
    .X(_0785_));
 sky130_fd_sc_hd__a221oi_1 _4069_ (.A1(_0458_),
    .A2(_0781_),
    .B1(_3037_),
    .B2(_0782_),
    .C1(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__clkbuf_4 _4070_ (.A(_3036_),
    .X(_0787_));
 sky130_fd_sc_hd__buf_4 _4071_ (.A(_3039_),
    .X(_0788_));
 sky130_fd_sc_hd__inv_2 _4072_ (.A(_2990_),
    .Y(_0789_));
 sky130_fd_sc_hd__clkbuf_4 _4073_ (.A(_3032_),
    .X(_0790_));
 sky130_fd_sc_hd__clkbuf_4 _4074_ (.A(_3033_),
    .X(_0791_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(_0791_),
    .B(_3030_),
    .Y(_0792_));
 sky130_fd_sc_hd__o21ai_1 _4076_ (.A1(_0789_),
    .A2(_0790_),
    .B1(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__a221oi_1 _4077_ (.A1(_3058_),
    .A2(_0787_),
    .B1(_0402_),
    .B2(_0788_),
    .C1(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _4078_ (.A(\egd_top.BitStream_buffer.BS_buffer[116] ),
    .Y(_0795_));
 sky130_fd_sc_hd__clkbuf_4 _4079_ (.A(_3068_),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_4 _4080_ (.A(_3069_),
    .X(_0797_));
 sky130_fd_sc_hd__nand2_1 _4081_ (.A(_0797_),
    .B(_2800_),
    .Y(_0798_));
 sky130_fd_sc_hd__o221a_1 _4082_ (.A1(_0795_),
    .A2(_3065_),
    .B1(_0723_),
    .B2(_0796_),
    .C1(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__clkbuf_4 _4083_ (.A(_3055_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_4 _4084_ (.A(_3056_),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_4 _4085_ (.A(_3057_),
    .X(_0802_));
 sky130_fd_sc_hd__nand2_1 _4086_ (.A(_0802_),
    .B(_3070_),
    .Y(_0803_));
 sky130_fd_sc_hd__clkbuf_4 _4087_ (.A(_3060_),
    .X(_0804_));
 sky130_fd_sc_hd__nand2_1 _4088_ (.A(_0804_),
    .B(_2820_),
    .Y(_0805_));
 sky130_fd_sc_hd__nand2_1 _4089_ (.A(_0803_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a221oi_1 _4090_ (.A1(_3066_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2812_),
    .C1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__and4_1 _4091_ (.A(_0786_),
    .B(_0794_),
    .C(_0799_),
    .D(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__clkbuf_4 _4092_ (.A(_2986_),
    .X(_0809_));
 sky130_fd_sc_hd__clkbuf_4 _4093_ (.A(_2989_),
    .X(_0810_));
 sky130_fd_sc_hd__buf_4 _4094_ (.A(_2982_),
    .X(_0811_));
 sky130_fd_sc_hd__clkbuf_4 _4095_ (.A(_2992_),
    .X(_0812_));
 sky130_fd_sc_hd__nand2_1 _4096_ (.A(_0812_),
    .B(_3040_),
    .Y(_0813_));
 sky130_fd_sc_hd__o21ai_1 _4097_ (.A1(_2908_),
    .A2(_0811_),
    .B1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a221oi_1 _4098_ (.A1(_3002_),
    .A2(_0809_),
    .B1(_3153_),
    .B2(_0810_),
    .C1(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__clkbuf_4 _4099_ (.A(_3001_),
    .X(_0816_));
 sky130_fd_sc_hd__clkbuf_4 _4100_ (.A(_2997_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _4101_ (.A(_2999_),
    .X(_0818_));
 sky130_fd_sc_hd__nand2_1 _4102_ (.A(_0818_),
    .B(_2816_),
    .Y(_0819_));
 sky130_fd_sc_hd__clkbuf_4 _4103_ (.A(_3004_),
    .X(_0820_));
 sky130_fd_sc_hd__nand2_1 _4104_ (.A(_0820_),
    .B(_2810_),
    .Y(_0821_));
 sky130_fd_sc_hd__nand2_1 _4105_ (.A(_0819_),
    .B(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__a221oi_1 _4106_ (.A1(_0816_),
    .A2(_3053_),
    .B1(_0817_),
    .B2(_2818_),
    .C1(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__clkbuf_4 _4107_ (.A(_3014_),
    .X(_0824_));
 sky130_fd_sc_hd__clkbuf_4 _4108_ (.A(_3016_),
    .X(_0825_));
 sky130_fd_sc_hd__clkbuf_4 _4109_ (.A(_3009_),
    .X(_0826_));
 sky130_fd_sc_hd__clkbuf_4 _4110_ (.A(_3012_),
    .X(_0827_));
 sky130_fd_sc_hd__o22ai_1 _4111_ (.A1(_0407_),
    .A2(_0826_),
    .B1(_0757_),
    .B2(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__a221oi_1 _4112_ (.A1(_0824_),
    .A2(_2863_),
    .B1(_0825_),
    .B2(_2920_),
    .C1(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__clkbuf_8 _4113_ (.A(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_4 _4114_ (.A(_3022_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_4 _4115_ (.A(_3020_),
    .X(_0832_));
 sky130_fd_sc_hd__clkbuf_4 _4116_ (.A(_3024_),
    .X(_0833_));
 sky130_fd_sc_hd__nand2_1 _4117_ (.A(_0833_),
    .B(_2808_),
    .Y(_0834_));
 sky130_fd_sc_hd__clkbuf_4 _4118_ (.A(_3026_),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _4119_ (.A(_0835_),
    .B(_2824_),
    .Y(_0836_));
 sky130_fd_sc_hd__nand2_1 _4120_ (.A(_0834_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__a221oi_1 _4121_ (.A1(_0830_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2814_),
    .C1(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__and4_1 _4122_ (.A(_0815_),
    .B(_0823_),
    .C(_0829_),
    .D(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__clkbuf_4 _4123_ (.A(_2896_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_8 _4124_ (.A(\egd_top.BitStream_buffer.BS_buffer[9] ),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_4 _4125_ (.A(_2900_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_4 _4126_ (.A(_2894_),
    .X(_0843_));
 sky130_fd_sc_hd__clkbuf_4 _4127_ (.A(_2903_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(_0844_),
    .B(_0610_),
    .Y(_0845_));
 sky130_fd_sc_hd__o21ai_1 _4129_ (.A1(_0546_),
    .A2(_0843_),
    .B1(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__a221oi_1 _4130_ (.A1(_0469_),
    .A2(_0840_),
    .B1(_0841_),
    .B2(_0842_),
    .C1(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__buf_4 _4131_ (.A(_2880_),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_4 _4132_ (.A(_2886_),
    .X(_0849_));
 sky130_fd_sc_hd__clkbuf_4 _4133_ (.A(_0629_),
    .X(_0850_));
 sky130_fd_sc_hd__nand2_1 _4134_ (.A(_2867_),
    .B(_2913_),
    .Y(_0851_));
 sky130_fd_sc_hd__o21ai_1 _4135_ (.A1(_0474_),
    .A2(_0850_),
    .B1(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__a221oi_1 _4136_ (.A1(_0414_),
    .A2(_0848_),
    .B1(_3010_),
    .B2(_0849_),
    .C1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _4137_ (.A(_2858_),
    .B(_2848_),
    .Y(_0854_));
 sky130_fd_sc_hd__o21ai_1 _4138_ (.A1(_0444_),
    .A2(_2854_),
    .B1(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__a221oi_1 _4139_ (.A1(_0464_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0495_),
    .C1(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__buf_4 _4140_ (.A(_2919_),
    .X(_0857_));
 sky130_fd_sc_hd__buf_4 _4141_ (.A(_2921_),
    .X(_0858_));
 sky130_fd_sc_hd__inv_2 _4142_ (.A(_0395_),
    .Y(_0859_));
 sky130_fd_sc_hd__o22ai_1 _4143_ (.A1(_0859_),
    .A2(_2912_),
    .B1(_3091_),
    .B2(_2917_),
    .Y(_0860_));
 sky130_fd_sc_hd__a221oi_1 _4144_ (.A1(_2980_),
    .A2(_0857_),
    .B1(_3097_),
    .B2(_0858_),
    .C1(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__and4_1 _4145_ (.A(_0847_),
    .B(_0853_),
    .C(_0856_),
    .D(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_8 _4146_ (.A(_2929_),
    .X(_0863_));
 sky130_fd_sc_hd__buf_4 _4147_ (.A(_2930_),
    .X(_0864_));
 sky130_fd_sc_hd__clkbuf_4 _4148_ (.A(_2934_),
    .X(_0865_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(_0865_),
    .B(_0343_),
    .Y(_0866_));
 sky130_fd_sc_hd__clkbuf_4 _4150_ (.A(_2938_),
    .X(_0867_));
 sky130_fd_sc_hd__nand2_1 _4151_ (.A(_0867_),
    .B(_3112_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand2_1 _4152_ (.A(_0866_),
    .B(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__a221oi_2 _4153_ (.A1(_3119_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_0346_),
    .C1(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__clkbuf_8 _4154_ (.A(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_0871_));
 sky130_fd_sc_hd__clkbuf_4 _4155_ (.A(_2976_),
    .X(_0872_));
 sky130_fd_sc_hd__clkbuf_4 _4156_ (.A(_2971_),
    .X(_0873_));
 sky130_fd_sc_hd__clkbuf_4 _4157_ (.A(_2969_),
    .X(_0874_));
 sky130_fd_sc_hd__clkbuf_8 _4158_ (.A(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .X(_0875_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(_0874_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__clkbuf_4 _4160_ (.A(_2973_),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _4161_ (.A(_0877_),
    .B(_0336_),
    .Y(_0878_));
 sky130_fd_sc_hd__nand2_1 _4162_ (.A(_0876_),
    .B(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__a221oi_1 _4163_ (.A1(_0871_),
    .A2(_0872_),
    .B1(_0657_),
    .B2(_0873_),
    .C1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__inv_2 _4164_ (.A(_2887_),
    .Y(_0881_));
 sky130_fd_sc_hd__buf_4 _4165_ (.A(_2945_),
    .X(_0882_));
 sky130_fd_sc_hd__clkbuf_4 _4166_ (.A(_2947_),
    .X(_0883_));
 sky130_fd_sc_hd__nand2_1 _4167_ (.A(_0883_),
    .B(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .Y(_0884_));
 sky130_fd_sc_hd__clkbuf_4 _4168_ (.A(_2949_),
    .X(_0885_));
 sky130_fd_sc_hd__clkbuf_8 _4169_ (.A(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .X(_0886_));
 sky130_fd_sc_hd__nand2_1 _4170_ (.A(_0885_),
    .B(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_2 _4171_ (.A(_3139_),
    .Y(_0888_));
 sky130_fd_sc_hd__buf_2 _4172_ (.A(_2953_),
    .X(_0889_));
 sky130_fd_sc_hd__or2_1 _4173_ (.A(_0888_),
    .B(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__o2111a_1 _4174_ (.A1(_0881_),
    .A2(_0882_),
    .B1(_0884_),
    .C1(_0887_),
    .D1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_4 _4175_ (.A(_2956_),
    .X(_0892_));
 sky130_fd_sc_hd__clkbuf_4 _4176_ (.A(_2958_),
    .X(_0893_));
 sky130_fd_sc_hd__buf_4 _4177_ (.A(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .X(_0894_));
 sky130_fd_sc_hd__clkbuf_4 _4178_ (.A(_2962_),
    .X(_0895_));
 sky130_fd_sc_hd__nand2_1 _4179_ (.A(_0895_),
    .B(\egd_top.BitStream_buffer.BS_buffer[124] ),
    .Y(_0896_));
 sky130_fd_sc_hd__clkbuf_4 _4180_ (.A(_2965_),
    .X(_0897_));
 sky130_fd_sc_hd__nand2_1 _4181_ (.A(_0897_),
    .B(_2830_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_1 _4182_ (.A(_0896_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__a221oi_1 _4183_ (.A1(_0892_),
    .A2(_3105_),
    .B1(_0893_),
    .B2(_0894_),
    .C1(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__and4_1 _4184_ (.A(_0870_),
    .B(_0880_),
    .C(_0891_),
    .D(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__and4_1 _4185_ (.A(_0808_),
    .B(_0839_),
    .C(_0862_),
    .D(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__buf_4 _4186_ (.A(_0456_),
    .X(_0903_));
 sky130_fd_sc_hd__inv_2 _4187_ (.A(_0385_),
    .Y(_0904_));
 sky130_fd_sc_hd__o22ai_1 _4188_ (.A1(_0904_),
    .A2(_3131_),
    .B1(_0731_),
    .B2(_3135_),
    .Y(_0905_));
 sky130_fd_sc_hd__a221oi_1 _4189_ (.A1(_2935_),
    .A2(_3126_),
    .B1(_0378_),
    .B2(_3123_),
    .C1(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__buf_4 _4190_ (.A(_3111_),
    .X(_0907_));
 sky130_fd_sc_hd__buf_4 _4191_ (.A(_3114_),
    .X(_0908_));
 sky130_fd_sc_hd__nand2_1 _4192_ (.A(_3118_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_0909_));
 sky130_fd_sc_hd__o21ai_1 _4193_ (.A1(_0717_),
    .A2(_3110_),
    .B1(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__a221oi_2 _4194_ (.A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .A2(_0907_),
    .B1(_2951_),
    .B2(_0908_),
    .C1(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _4195_ (.A(_3100_),
    .B(_2943_),
    .Y(_0912_));
 sky130_fd_sc_hd__o21ai_1 _4196_ (.A1(_0641_),
    .A2(_3093_),
    .B1(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__a221oi_1 _4197_ (.A1(_3127_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_2859_),
    .C1(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__or2_1 _4198_ (.A(_0489_),
    .B(_3080_),
    .X(_0915_));
 sky130_fd_sc_hd__or2_1 _4199_ (.A(_0544_),
    .B(_3084_),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _4200_ (.A(_3087_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_0917_));
 sky130_fd_sc_hd__o2111a_1 _4201_ (.A1(_3129_),
    .A2(_3077_),
    .B1(_0915_),
    .C1(_0916_),
    .D1(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__and4_1 _4202_ (.A(_0906_),
    .B(_0911_),
    .C(_0914_),
    .D(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_8 _4203_ (.A(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_4 _4204_ (.A(_0361_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_4 _4205_ (.A(_0363_),
    .X(_0922_));
 sky130_fd_sc_hd__buf_4 _4206_ (.A(_0357_),
    .X(_0923_));
 sky130_fd_sc_hd__or2b_1 _4207_ (.A(_0923_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_4 _4208_ (.A(_0359_),
    .X(_0925_));
 sky130_fd_sc_hd__buf_4 _4209_ (.A(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .X(_0926_));
 sky130_fd_sc_hd__nand2_1 _4210_ (.A(_0925_),
    .B(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__nand2_1 _4211_ (.A(_0924_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__a221oi_1 _4212_ (.A1(_0920_),
    .A2(_0921_),
    .B1(_0420_),
    .B2(_0922_),
    .C1(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__clkbuf_4 _4213_ (.A(_0368_),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_4 _4214_ (.A(_0370_),
    .X(_0931_));
 sky130_fd_sc_hd__a22o_1 _4215_ (.A1(_0371_),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_0553_),
    .X(_0932_));
 sky130_fd_sc_hd__clkbuf_4 _4216_ (.A(_0373_),
    .X(_0933_));
 sky130_fd_sc_hd__clkbuf_4 _4217_ (.A(_0374_),
    .X(_0934_));
 sky130_fd_sc_hd__a22o_1 _4218_ (.A1(_0933_),
    .A2(_0742_),
    .B1(_0934_),
    .B2(_0583_),
    .X(_0935_));
 sky130_fd_sc_hd__nor2_1 _4219_ (.A(_0932_),
    .B(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__clkbuf_4 _4220_ (.A(_0388_),
    .X(_0937_));
 sky130_fd_sc_hd__buf_4 _4221_ (.A(_0391_),
    .X(_0938_));
 sky130_fd_sc_hd__clkbuf_4 _4222_ (.A(_0394_),
    .X(_0939_));
 sky130_fd_sc_hd__nand2_1 _4223_ (.A(_0939_),
    .B(_0341_),
    .Y(_0940_));
 sky130_fd_sc_hd__clkbuf_4 _4224_ (.A(_0397_),
    .X(_0941_));
 sky130_fd_sc_hd__nand2_1 _4225_ (.A(_0941_),
    .B(_2957_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _4226_ (.A(_0940_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__a221oi_2 _4227_ (.A1(_0937_),
    .A2(_3142_),
    .B1(_0398_),
    .B2(_0938_),
    .C1(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__clkbuf_4 _4228_ (.A(_0380_),
    .X(_0945_));
 sky130_fd_sc_hd__buf_4 _4229_ (.A(_0377_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_4 _4230_ (.A(_0382_),
    .X(_0947_));
 sky130_fd_sc_hd__nand2_1 _4231_ (.A(_0947_),
    .B(_0389_),
    .Y(_0948_));
 sky130_fd_sc_hd__clkbuf_4 _4232_ (.A(_0384_),
    .X(_0949_));
 sky130_fd_sc_hd__nand2_1 _4233_ (.A(_0949_),
    .B(_0392_),
    .Y(_0950_));
 sky130_fd_sc_hd__nand2_1 _4234_ (.A(_0948_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__a221oi_1 _4235_ (.A1(_0463_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_2974_),
    .C1(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__and4_2 _4236_ (.A(_0929_),
    .B(_0936_),
    .C(_0944_),
    .D(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__buf_6 _4237_ (.A(_3157_),
    .X(_0954_));
 sky130_fd_sc_hd__buf_8 _4238_ (.A(_0329_),
    .X(_0955_));
 sky130_fd_sc_hd__buf_4 _4239_ (.A(_3152_),
    .X(_0956_));
 sky130_fd_sc_hd__inv_2 _4240_ (.A(\egd_top.BitStream_buffer.BS_buffer[112] ),
    .Y(_0957_));
 sky130_fd_sc_hd__buf_4 _4241_ (.A(_3155_),
    .X(_0958_));
 sky130_fd_sc_hd__o22ai_1 _4242_ (.A1(_0772_),
    .A2(_0956_),
    .B1(_0957_),
    .B2(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__a221oi_2 _4243_ (.A1(_2804_),
    .A2(_0954_),
    .B1(_2802_),
    .B2(_0955_),
    .C1(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__clkbuf_4 _4244_ (.A(_3141_),
    .X(_0961_));
 sky130_fd_sc_hd__clkbuf_4 _4245_ (.A(_2771_),
    .X(_0962_));
 sky130_fd_sc_hd__clkbuf_4 _4246_ (.A(_3145_),
    .X(_0963_));
 sky130_fd_sc_hd__clkbuf_4 _4247_ (.A(_3148_),
    .X(_0964_));
 sky130_fd_sc_hd__o22ai_1 _4248_ (.A1(_3133_),
    .A2(_0963_),
    .B1(_0575_),
    .B2(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__a221oi_1 _4249_ (.A1(_0435_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_0366_),
    .C1(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__clkbuf_4 _4250_ (.A(_0352_),
    .X(_0967_));
 sky130_fd_sc_hd__clkbuf_4 _4251_ (.A(_0353_),
    .X(_0968_));
 sky130_fd_sc_hd__clkbuf_4 _4252_ (.A(_0348_),
    .X(_0969_));
 sky130_fd_sc_hd__inv_2 _4253_ (.A(_2926_),
    .Y(_0970_));
 sky130_fd_sc_hd__clkbuf_4 _4254_ (.A(_0350_),
    .X(_0971_));
 sky130_fd_sc_hd__o22ai_1 _4255_ (.A1(_3075_),
    .A2(_0969_),
    .B1(_0970_),
    .B2(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__a221oi_1 _4256_ (.A1(_0967_),
    .A2(_0625_),
    .B1(_0968_),
    .B2(_0777_),
    .C1(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__clkbuf_4 _4257_ (.A(_0340_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_4 _4258_ (.A(_0342_),
    .X(_0975_));
 sky130_fd_sc_hd__clkbuf_4 _4259_ (.A(_0335_),
    .X(_0976_));
 sky130_fd_sc_hd__clkbuf_4 _4260_ (.A(_0338_),
    .X(_0977_));
 sky130_fd_sc_hd__o22ai_1 _4261_ (.A1(_3147_),
    .A2(_0976_),
    .B1(_0349_),
    .B2(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__a221oi_1 _4262_ (.A1(_0974_),
    .A2(_0333_),
    .B1(_0975_),
    .B2(_3143_),
    .C1(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__and4_1 _4263_ (.A(_0960_),
    .B(_0966_),
    .C(_0973_),
    .D(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_4 _4264_ (.A(_0411_),
    .X(_0981_));
 sky130_fd_sc_hd__clkbuf_4 _4265_ (.A(_0413_),
    .X(_0982_));
 sky130_fd_sc_hd__inv_2 _4266_ (.A(_2922_),
    .Y(_0983_));
 sky130_fd_sc_hd__inv_2 _4267_ (.A(_3017_),
    .Y(_0984_));
 sky130_fd_sc_hd__o22ai_1 _4268_ (.A1(_0983_),
    .A2(_0405_),
    .B1(_0984_),
    .B2(_0409_),
    .Y(_0985_));
 sky130_fd_sc_hd__a221oi_1 _4269_ (.A1(_0981_),
    .A2(_3007_),
    .B1(_0982_),
    .B2(_2993_),
    .C1(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__buf_4 _4270_ (.A(_0422_),
    .X(_0987_));
 sky130_fd_sc_hd__buf_6 _4271_ (.A(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .X(_0988_));
 sky130_fd_sc_hd__buf_4 _4272_ (.A(_0417_),
    .X(_0989_));
 sky130_fd_sc_hd__buf_4 _4273_ (.A(_0419_),
    .X(_0990_));
 sky130_fd_sc_hd__nand2_1 _4274_ (.A(_0990_),
    .B(_0477_),
    .Y(_0991_));
 sky130_fd_sc_hd__clkbuf_4 _4275_ (.A(_0424_),
    .X(_0992_));
 sky130_fd_sc_hd__nand2_1 _4276_ (.A(_0992_),
    .B(_2987_),
    .Y(_0993_));
 sky130_fd_sc_hd__nand2_1 _4277_ (.A(_0991_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__a221oi_2 _4278_ (.A1(_0551_),
    .A2(_0987_),
    .B1(_0988_),
    .B2(_0989_),
    .C1(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__clkbuf_4 _4279_ (.A(_0434_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_4 _4280_ (.A(_0430_),
    .X(_0997_));
 sky130_fd_sc_hd__nand2_1 _4281_ (.A(_0428_),
    .B(_2959_),
    .Y(_0998_));
 sky130_fd_sc_hd__clkbuf_4 _4282_ (.A(_0432_),
    .X(_0999_));
 sky130_fd_sc_hd__buf_4 _4283_ (.A(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .X(_1000_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_0999_),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_0998_),
    .B(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__a221oi_1 _4286_ (.A1(_0656_),
    .A2(_0996_),
    .B1(_0709_),
    .B2(_0997_),
    .C1(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__a22o_1 _4287_ (.A1(_0439_),
    .A2(_0607_),
    .B1(_0441_),
    .B2(_2904_),
    .X(_1004_));
 sky130_fd_sc_hd__inv_2 _4288_ (.A(\egd_top.BitStream_buffer.BS_buffer[101] ),
    .Y(_1005_));
 sky130_fd_sc_hd__o22ai_1 _4289_ (.A1(_1005_),
    .A2(_0446_),
    .B1(_0465_),
    .B2(_0449_),
    .Y(_1006_));
 sky130_fd_sc_hd__nor2_1 _4290_ (.A(_1004_),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__and4_1 _4291_ (.A(_0986_),
    .B(_0995_),
    .C(_1003_),
    .D(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__and4_1 _4292_ (.A(_0919_),
    .B(_0953_),
    .C(_0980_),
    .D(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nand3_1 _4293_ (.A(_0902_),
    .B(_0903_),
    .C(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__clkbuf_8 _4294_ (.A(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .X(_1011_));
 sky130_fd_sc_hd__o21a_1 _4295_ (.A1(_1011_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1012_));
 sky130_fd_sc_hd__nand2_1 _4296_ (.A(_1010_),
    .B(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__nand2_1 _4297_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_1014_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_1013_),
    .B(_1014_),
    .Y(_0301_));
 sky130_fd_sc_hd__a22o_1 _4299_ (.A1(\egd_top.BitStream_buffer.BS_buffer[127] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0458_),
    .X(_1015_));
 sky130_fd_sc_hd__a221oi_1 _4300_ (.A1(_0625_),
    .A2(_0781_),
    .B1(_3053_),
    .B2(_0782_),
    .C1(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__clkinv_4 _4301_ (.A(_3058_),
    .Y(_1017_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_0791_),
    .B(_3037_),
    .Y(_1018_));
 sky130_fd_sc_hd__o21ai_1 _4303_ (.A1(_1017_),
    .A2(_0790_),
    .B1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__a221oi_1 _4304_ (.A1(_3066_),
    .A2(_0787_),
    .B1(_2863_),
    .B2(_0788_),
    .C1(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__inv_2 _4305_ (.A(\egd_top.BitStream_buffer.BS_buffer[117] ),
    .Y(_1021_));
 sky130_fd_sc_hd__nand2_1 _4306_ (.A(_0797_),
    .B(_2802_),
    .Y(_1022_));
 sky130_fd_sc_hd__o221a_1 _4307_ (.A1(_1021_),
    .A2(_3065_),
    .B1(_0957_),
    .B2(_0796_),
    .C1(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__nand2_1 _4308_ (.A(_0802_),
    .B(_0330_),
    .Y(_1024_));
 sky130_fd_sc_hd__nand2_1 _4309_ (.A(_0804_),
    .B(_2822_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(_1024_),
    .B(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__a221oi_1 _4311_ (.A1(_3153_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2814_),
    .C1(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__and4_1 _4312_ (.A(_1016_),
    .B(_1020_),
    .C(_1023_),
    .D(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__nand2_1 _4313_ (.A(_0812_),
    .B(_3015_),
    .Y(_1029_));
 sky130_fd_sc_hd__o21ai_1 _4314_ (.A1(_0480_),
    .A2(_0811_),
    .B1(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__a221oi_1 _4315_ (.A1(_3030_),
    .A2(_0809_),
    .B1(_3070_),
    .B2(_0810_),
    .C1(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__nand2_1 _4316_ (.A(_0818_),
    .B(_2818_),
    .Y(_1032_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_0820_),
    .B(_2812_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(_1032_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__a221oi_1 _4319_ (.A1(_0816_),
    .A2(_2990_),
    .B1(_0817_),
    .B2(_2820_),
    .C1(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__o22ai_1 _4320_ (.A1(_0602_),
    .A2(_0826_),
    .B1(_0984_),
    .B2(_0827_),
    .Y(_1036_));
 sky130_fd_sc_hd__a221oi_1 _4321_ (.A1(_0824_),
    .A2(_2920_),
    .B1(_0825_),
    .B2(_2922_),
    .C1(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(_0833_),
    .B(_2810_),
    .Y(_1038_));
 sky130_fd_sc_hd__nand2_1 _4323_ (.A(_0835_),
    .B(_2826_),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _4324_ (.A(_1038_),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__a221oi_1 _4325_ (.A1(_0926_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2816_),
    .C1(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__and4_1 _4326_ (.A(_1031_),
    .B(_1035_),
    .C(_1037_),
    .D(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__nand2_1 _4327_ (.A(_0844_),
    .B(_0443_),
    .Y(_1043_));
 sky130_fd_sc_hd__o21ai_1 _4328_ (.A1(_3078_),
    .A2(_0843_),
    .B1(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__a221oi_1 _4329_ (.A1(_0988_),
    .A2(_0840_),
    .B1(_3101_),
    .B2(_0842_),
    .C1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__nand2_1 _4330_ (.A(_2867_),
    .B(_2980_),
    .Y(_1046_));
 sky130_fd_sc_hd__o21ai_1 _4331_ (.A1(_3082_),
    .A2(_0850_),
    .B1(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__a221oi_1 _4332_ (.A1(_2887_),
    .A2(_0848_),
    .B1(_0406_),
    .B2(_0849_),
    .C1(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(_2858_),
    .B(_0464_),
    .Y(_1049_));
 sky130_fd_sc_hd__o21ai_1 _4334_ (.A1(_0619_),
    .A2(_2854_),
    .B1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__a221oi_2 _4335_ (.A1(_2959_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0657_),
    .C1(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__inv_2 _4336_ (.A(_2935_),
    .Y(_1052_));
 sky130_fd_sc_hd__o22ai_1 _4337_ (.A1(_1052_),
    .A2(_2912_),
    .B1(_2908_),
    .B2(_2917_),
    .Y(_1053_));
 sky130_fd_sc_hd__a221oi_1 _4338_ (.A1(_3097_),
    .A2(_0857_),
    .B1(_3090_),
    .B2(_0858_),
    .C1(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__and4_1 _4339_ (.A(_1045_),
    .B(_1048_),
    .C(_1051_),
    .D(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_1 _4340_ (.A(_0865_),
    .B(_2974_),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_1 _4341_ (.A(_0867_),
    .B(_3119_),
    .Y(_1057_));
 sky130_fd_sc_hd__nand2_1 _4342_ (.A(_1056_),
    .B(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__a221oi_2 _4343_ (.A1(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_3112_),
    .C1(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__nand2_1 _4344_ (.A(_0874_),
    .B(_0587_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand2_1 _4345_ (.A(_0877_),
    .B(_3146_),
    .Y(_1061_));
 sky130_fd_sc_hd__nand2_1 _4346_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a221oi_1 _4347_ (.A1(_0420_),
    .A2(_0872_),
    .B1(_0894_),
    .B2(_0873_),
    .C1(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__nand2_1 _4348_ (.A(_0883_),
    .B(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .Y(_1064_));
 sky130_fd_sc_hd__nand2_1 _4349_ (.A(_0885_),
    .B(_2874_),
    .Y(_1065_));
 sky130_fd_sc_hd__inv_2 _4350_ (.A(\egd_top.BitStream_buffer.BS_buffer[65] ),
    .Y(_1066_));
 sky130_fd_sc_hd__or2_1 _4351_ (.A(_1066_),
    .B(_0889_),
    .X(_1067_));
 sky130_fd_sc_hd__o2111a_1 _4352_ (.A1(_3008_),
    .A2(_0882_),
    .B1(_1064_),
    .C1(_1065_),
    .D1(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__nand2_1 _4353_ (.A(_0895_),
    .B(\egd_top.BitStream_buffer.BS_buffer[125] ),
    .Y(_1069_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_0897_),
    .B(_0463_),
    .Y(_1070_));
 sky130_fd_sc_hd__nand2_1 _4355_ (.A(_1069_),
    .B(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__a221oi_1 _4356_ (.A1(_0892_),
    .A2(_0553_),
    .B1(_0893_),
    .B2(_1000_),
    .C1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__and4_1 _4357_ (.A(_1059_),
    .B(_1063_),
    .C(_1068_),
    .D(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__and4_1 _4358_ (.A(_1028_),
    .B(_1042_),
    .C(_1055_),
    .D(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__inv_2 _4359_ (.A(_0389_),
    .Y(_1075_));
 sky130_fd_sc_hd__o22ai_1 _4360_ (.A1(_1075_),
    .A2(_3131_),
    .B1(_0970_),
    .B2(_3135_),
    .Y(_1076_));
 sky130_fd_sc_hd__a221oi_2 _4361_ (.A1(_0378_),
    .A2(_3126_),
    .B1(_0341_),
    .B2(_3123_),
    .C1(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__nand2_1 _4362_ (.A(_3118_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1078_));
 sky130_fd_sc_hd__o21ai_1 _4363_ (.A1(_0904_),
    .A2(_3110_),
    .B1(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__a221oi_1 _4364_ (.A1(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .A2(_0907_),
    .B1(_0392_),
    .B2(_0908_),
    .C1(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(_3100_),
    .B(_0412_),
    .Y(_1081_));
 sky130_fd_sc_hd__o21ai_1 _4366_ (.A1(_0859_),
    .A2(_3093_),
    .B1(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__a221oi_2 _4367_ (.A1(_3124_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_2830_),
    .C1(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__or2_1 _4368_ (.A(_0650_),
    .B(_3080_),
    .X(_1084_));
 sky130_fd_sc_hd__or2_1 _4369_ (.A(_2944_),
    .B(_3084_),
    .X(_1085_));
 sky130_fd_sc_hd__nand2_1 _4370_ (.A(_3087_),
    .B(_3115_),
    .Y(_1086_));
 sky130_fd_sc_hd__o2111a_1 _4371_ (.A1(_0561_),
    .A2(_3077_),
    .B1(_1084_),
    .C1(_1085_),
    .D1(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__and4_1 _4372_ (.A(_1077_),
    .B(_1080_),
    .C(_1083_),
    .D(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__or2b_1 _4373_ (.A(_0923_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .X(_1089_));
 sky130_fd_sc_hd__nand2_1 _4374_ (.A(_0925_),
    .B(_0920_),
    .Y(_1090_));
 sky130_fd_sc_hd__nand2_1 _4375_ (.A(_1089_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__a221oi_1 _4376_ (.A1(_0875_),
    .A2(_0921_),
    .B1(_0607_),
    .B2(_0922_),
    .C1(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__a22o_1 _4377_ (.A1(_0656_),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_0709_),
    .X(_1093_));
 sky130_fd_sc_hd__a22o_1 _4378_ (.A1(_0933_),
    .A2(_0583_),
    .B1(_0934_),
    .B2(_0871_),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_1 _4379_ (.A(_1093_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(_0939_),
    .B(_0343_),
    .Y(_1096_));
 sky130_fd_sc_hd__nand2_1 _4381_ (.A(_0941_),
    .B(_0371_),
    .Y(_1097_));
 sky130_fd_sc_hd__nand2_1 _4382_ (.A(_1096_),
    .B(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__a221oi_1 _4383_ (.A1(_0937_),
    .A2(_3139_),
    .B1(_0366_),
    .B2(_0938_),
    .C1(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__nand2_1 _4384_ (.A(_0947_),
    .B(_2951_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _4385_ (.A(_0949_),
    .B(_3142_),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2_1 _4386_ (.A(_1100_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__a221oi_1 _4387_ (.A1(_2848_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_0333_),
    .C1(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__and4_1 _4388_ (.A(_1092_),
    .B(_1095_),
    .C(_1099_),
    .D(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__o22ai_2 _4389_ (.A1(_1005_),
    .A2(_0956_),
    .B1(_3064_),
    .B2(_0958_),
    .Y(_1105_));
 sky130_fd_sc_hd__a221oi_2 _4390_ (.A1(_2806_),
    .A2(_0954_),
    .B1(_2804_),
    .B2(_0955_),
    .C1(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__o22ai_1 _4391_ (.A1(_0349_),
    .A2(_0963_),
    .B1(_0731_),
    .B2(_0964_),
    .Y(_1107_));
 sky130_fd_sc_hd__a221oi_1 _4392_ (.A1(_2957_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_0435_),
    .C1(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__o22ai_1 _4393_ (.A1(_0543_),
    .A2(_0969_),
    .B1(_0347_),
    .B2(_0971_),
    .Y(_1109_));
 sky130_fd_sc_hd__a221oi_1 _4394_ (.A1(_0967_),
    .A2(_0777_),
    .B1(_0968_),
    .B2(_1011_),
    .C1(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__o22ai_1 _4395_ (.A1(_3133_),
    .A2(_0976_),
    .B1(_0575_),
    .B2(_0977_),
    .Y(_1111_));
 sky130_fd_sc_hd__a221oi_1 _4396_ (.A1(_0974_),
    .A2(_3143_),
    .B1(_0975_),
    .B2(_0336_),
    .C1(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__and4_1 _4397_ (.A(_1106_),
    .B(_1108_),
    .C(_1110_),
    .D(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__o22ai_1 _4398_ (.A1(_2914_),
    .A2(_0405_),
    .B1(_0403_),
    .B2(_0409_),
    .Y(_1114_));
 sky130_fd_sc_hd__a221oi_1 _4399_ (.A1(_0981_),
    .A2(_2993_),
    .B1(_0982_),
    .B2(_3010_),
    .C1(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__clkbuf_8 _4400_ (.A(\egd_top.BitStream_buffer.BS_buffer[8] ),
    .X(_1116_));
 sky130_fd_sc_hd__nand2_1 _4401_ (.A(_0990_),
    .B(_0638_),
    .Y(_1117_));
 sky130_fd_sc_hd__nand2_1 _4402_ (.A(_0992_),
    .B(_3034_),
    .Y(_1118_));
 sky130_fd_sc_hd__nand2_1 _4403_ (.A(_1117_),
    .B(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__a221oi_2 _4404_ (.A1(_2881_),
    .A2(_0987_),
    .B1(_1116_),
    .B2(_0989_),
    .C1(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(_0428_),
    .B(_0495_),
    .Y(_1121_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_0999_),
    .B(_0830_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand2_1 _4407_ (.A(_1121_),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__a221oi_1 _4408_ (.A1(_3105_),
    .A2(_0996_),
    .B1(_2859_),
    .B2(_0997_),
    .C1(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__a22o_1 _4409_ (.A1(_0439_),
    .A2(_2904_),
    .B1(_0441_),
    .B2(_0477_),
    .X(_1125_));
 sky130_fd_sc_hd__clkinv_4 _4410_ (.A(\egd_top.BitStream_buffer.BS_buffer[102] ),
    .Y(_1126_));
 sky130_fd_sc_hd__o22ai_1 _4411_ (.A1(_1126_),
    .A2(_0446_),
    .B1(_3151_),
    .B2(_0449_),
    .Y(_1127_));
 sky130_fd_sc_hd__nor2_1 _4412_ (.A(_1125_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__and4_1 _4413_ (.A(_1115_),
    .B(_1120_),
    .C(_1124_),
    .D(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__and4_1 _4414_ (.A(_1088_),
    .B(_1104_),
    .C(_1113_),
    .D(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__nand3_1 _4415_ (.A(_1074_),
    .B(_0903_),
    .C(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__o21a_1 _4416_ (.A1(_0886_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1132_));
 sky130_fd_sc_hd__nand2_1 _4417_ (.A(_1131_),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__nand2_1 _4418_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_1134_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_1133_),
    .B(_1134_),
    .Y(_0300_));
 sky130_fd_sc_hd__a22o_1 _4420_ (.A1(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0625_),
    .X(_1135_));
 sky130_fd_sc_hd__a221oi_1 _4421_ (.A1(_0777_),
    .A2(_0781_),
    .B1(_2990_),
    .B2(_0782_),
    .C1(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__nand2_1 _4422_ (.A(_0791_),
    .B(_3053_),
    .Y(_1137_));
 sky130_fd_sc_hd__o21ai_1 _4423_ (.A1(_3067_),
    .A2(_0790_),
    .B1(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__a221oi_1 _4424_ (.A1(_3153_),
    .A2(_0787_),
    .B1(_2920_),
    .B2(_0788_),
    .C1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__inv_2 _4425_ (.A(\egd_top.BitStream_buffer.BS_buffer[118] ),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _4426_ (.A(_0797_),
    .B(_2804_),
    .Y(_1141_));
 sky130_fd_sc_hd__o221a_1 _4427_ (.A1(_1140_),
    .A2(_3065_),
    .B1(_3064_),
    .B2(_0796_),
    .C1(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(_0802_),
    .B(_2791_),
    .Y(_1143_));
 sky130_fd_sc_hd__nand2_1 _4429_ (.A(_0804_),
    .B(_2824_),
    .Y(_1144_));
 sky130_fd_sc_hd__nand2_1 _4430_ (.A(_1143_),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__a221oi_1 _4431_ (.A1(_3070_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2816_),
    .C1(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__and4_1 _4432_ (.A(_1136_),
    .B(_1139_),
    .C(_1142_),
    .D(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nand2_1 _4433_ (.A(_0812_),
    .B(_3017_),
    .Y(_1148_));
 sky130_fd_sc_hd__o21ai_1 _4434_ (.A1(_0641_),
    .A2(_0811_),
    .B1(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__a221oi_1 _4435_ (.A1(_3037_),
    .A2(_0809_),
    .B1(_0330_),
    .B2(_0810_),
    .C1(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_1 _4436_ (.A(_0818_),
    .B(_2820_),
    .Y(_1151_));
 sky130_fd_sc_hd__nand2_1 _4437_ (.A(_0820_),
    .B(_2814_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(_1151_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__a221oi_1 _4439_ (.A1(_0816_),
    .A2(_3058_),
    .B1(_0817_),
    .B2(_2822_),
    .C1(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__o22ai_1 _4440_ (.A1(_0757_),
    .A2(_0826_),
    .B1(_0403_),
    .B2(_0827_),
    .Y(_1155_));
 sky130_fd_sc_hd__a221oi_1 _4441_ (.A1(_0824_),
    .A2(_2922_),
    .B1(_0825_),
    .B2(_2913_),
    .C1(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(_0833_),
    .B(_2812_),
    .Y(_1157_));
 sky130_fd_sc_hd__nand2_1 _4443_ (.A(_0835_),
    .B(_2828_),
    .Y(_1158_));
 sky130_fd_sc_hd__nand2_1 _4444_ (.A(_1157_),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__a221oi_2 _4445_ (.A1(_0920_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2818_),
    .C1(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__and4_1 _4446_ (.A(_1150_),
    .B(_1154_),
    .C(_1156_),
    .D(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(_0844_),
    .B(_2987_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21ai_1 _4448_ (.A1(_0544_),
    .A2(_0843_),
    .B1(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__a221oi_1 _4449_ (.A1(_1116_),
    .A2(_0840_),
    .B1(_0551_),
    .B2(_0842_),
    .C1(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__nand2_1 _4450_ (.A(_2867_),
    .B(_3097_),
    .Y(_1165_));
 sky130_fd_sc_hd__o21ai_1 _4451_ (.A1(_0546_),
    .A2(_0850_),
    .B1(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__a221oi_1 _4452_ (.A1(_3007_),
    .A2(_0848_),
    .B1(_3040_),
    .B2(_0849_),
    .C1(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__nand2_1 _4453_ (.A(_2858_),
    .B(_2959_),
    .Y(_1168_));
 sky130_fd_sc_hd__o21ai_1 _4454_ (.A1(_0772_),
    .A2(_2854_),
    .B1(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hd__a221oi_1 _4455_ (.A1(_0495_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0894_),
    .C1(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__inv_2 _4456_ (.A(_0378_),
    .Y(_1171_));
 sky130_fd_sc_hd__o22ai_1 _4457_ (.A1(_1171_),
    .A2(_2912_),
    .B1(_0480_),
    .B2(_2917_),
    .Y(_1172_));
 sky130_fd_sc_hd__a221oi_1 _4458_ (.A1(_3090_),
    .A2(_0857_),
    .B1(_2907_),
    .B2(_0858_),
    .C1(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__and4_1 _4459_ (.A(_1164_),
    .B(_1167_),
    .C(_1170_),
    .D(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_0865_),
    .B(_0333_),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_0867_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_1176_));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(_1175_),
    .B(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__a221oi_2 _4463_ (.A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_3119_),
    .C1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__nand2_1 _4464_ (.A(_0874_),
    .B(_0742_),
    .Y(_1179_));
 sky130_fd_sc_hd__nand2_1 _4465_ (.A(_0877_),
    .B(_3132_),
    .Y(_1180_));
 sky130_fd_sc_hd__nand2_1 _4466_ (.A(_1179_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__a221oi_1 _4467_ (.A1(_0607_),
    .A2(_0872_),
    .B1(_1000_),
    .B2(_0873_),
    .C1(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hd__nand2_1 _4468_ (.A(_0883_),
    .B(\egd_top.BitStream_buffer.BS_buffer[7] ),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _4469_ (.A(_0885_),
    .B(_0469_),
    .Y(_1184_));
 sky130_fd_sc_hd__inv_2 _4470_ (.A(\egd_top.BitStream_buffer.BS_buffer[66] ),
    .Y(_1185_));
 sky130_fd_sc_hd__or2_1 _4471_ (.A(_1185_),
    .B(_0889_),
    .X(_1186_));
 sky130_fd_sc_hd__o2111a_1 _4472_ (.A1(_0516_),
    .A2(_0882_),
    .B1(_1183_),
    .C1(_1184_),
    .D1(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__nand2_1 _4473_ (.A(_0895_),
    .B(_2826_),
    .Y(_1188_));
 sky130_fd_sc_hd__nand2_1 _4474_ (.A(_0897_),
    .B(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _4475_ (.A(_1188_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__a221oi_1 _4476_ (.A1(_0892_),
    .A2(_0709_),
    .B1(_0893_),
    .B2(_0830_),
    .C1(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__and4_1 _4477_ (.A(_1178_),
    .B(_1182_),
    .C(_1187_),
    .D(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__and4_1 _4478_ (.A(_1147_),
    .B(_1161_),
    .C(_1174_),
    .D(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__o22ai_1 _4479_ (.A1(_2952_),
    .A2(_3131_),
    .B1(_0347_),
    .B2(_3135_),
    .Y(_1194_));
 sky130_fd_sc_hd__a221oi_1 _4480_ (.A1(_0341_),
    .A2(_3126_),
    .B1(_0343_),
    .B2(_3123_),
    .C1(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_3118_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_1196_));
 sky130_fd_sc_hd__o21ai_1 _4482_ (.A1(_1075_),
    .A2(_3110_),
    .B1(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__a221oi_1 _4483_ (.A1(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .A2(_0907_),
    .B1(_3142_),
    .B2(_0908_),
    .C1(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__nand2_1 _4484_ (.A(_3100_),
    .B(_0414_),
    .Y(_1199_));
 sky130_fd_sc_hd__o21ai_1 _4485_ (.A1(_1052_),
    .A2(_3093_),
    .B1(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__a221oi_1 _4486_ (.A1(_0395_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_0463_),
    .C1(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__or2_1 _4487_ (.A(_0881_),
    .B(_3080_),
    .X(_1202_));
 sky130_fd_sc_hd__or2_1 _4488_ (.A(_0489_),
    .B(_3084_),
    .X(_1203_));
 sky130_fd_sc_hd__nand2_1 _4489_ (.A(_3087_),
    .B(_0385_),
    .Y(_1204_));
 sky130_fd_sc_hd__o2111a_1 _4490_ (.A1(_0717_),
    .A2(_3077_),
    .B1(_1202_),
    .C1(_1203_),
    .D1(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__and4_1 _4491_ (.A(_1195_),
    .B(_1198_),
    .C(_1201_),
    .D(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__or2b_1 _4492_ (.A(_0923_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .X(_1207_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(_0925_),
    .B(_0875_),
    .Y(_1208_));
 sky130_fd_sc_hd__nand2_1 _4494_ (.A(_1207_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__a221oi_1 _4495_ (.A1(_0587_),
    .A2(_0921_),
    .B1(_2904_),
    .B2(_0922_),
    .C1(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__a22o_1 _4496_ (.A1(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_2859_),
    .X(_1211_));
 sky130_fd_sc_hd__a22o_1 _4497_ (.A1(_0933_),
    .A2(_0871_),
    .B1(_0934_),
    .B2(_0420_),
    .X(_1212_));
 sky130_fd_sc_hd__nor2_1 _4498_ (.A(_1211_),
    .B(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_0939_),
    .B(_2974_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _4500_ (.A(_0941_),
    .B(_0656_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_1 _4501_ (.A(_1214_),
    .B(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__a221oi_1 _4502_ (.A1(_0937_),
    .A2(_0398_),
    .B1(_0435_),
    .B2(_0938_),
    .C1(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__nand2_1 _4503_ (.A(_0947_),
    .B(_0392_),
    .Y(_1218_));
 sky130_fd_sc_hd__nand2_1 _4504_ (.A(_0949_),
    .B(_3139_),
    .Y(_1219_));
 sky130_fd_sc_hd__nand2_1 _4505_ (.A(_1218_),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__a221oi_1 _4506_ (.A1(_0464_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_3143_),
    .C1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__and4_2 _4507_ (.A(_1210_),
    .B(_1213_),
    .C(_1217_),
    .D(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__o22ai_1 _4508_ (.A1(_1126_),
    .A2(_0956_),
    .B1(_0538_),
    .B2(_0958_),
    .Y(_1223_));
 sky130_fd_sc_hd__a221oi_2 _4509_ (.A1(_2808_),
    .A2(_0954_),
    .B1(_2806_),
    .B2(_0955_),
    .C1(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__o22ai_1 _4510_ (.A1(_0575_),
    .A2(_0963_),
    .B1(_0970_),
    .B2(_0964_),
    .Y(_1225_));
 sky130_fd_sc_hd__a221oi_1 _4511_ (.A1(_0371_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_2957_),
    .C1(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__o22ai_1 _4512_ (.A1(_3108_),
    .A2(_0969_),
    .B1(_0574_),
    .B2(_0971_),
    .Y(_1227_));
 sky130_fd_sc_hd__a221oi_1 _4513_ (.A1(_0967_),
    .A2(_1011_),
    .B1(_0968_),
    .B2(_0886_),
    .C1(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__o22ai_1 _4514_ (.A1(_0349_),
    .A2(_0976_),
    .B1(_0731_),
    .B2(_0977_),
    .Y(_1229_));
 sky130_fd_sc_hd__a221oi_1 _4515_ (.A1(_0974_),
    .A2(_0336_),
    .B1(_0975_),
    .B2(_3146_),
    .C1(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__and4_1 _4516_ (.A(_1224_),
    .B(_1226_),
    .C(_1228_),
    .D(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__o22ai_1 _4517_ (.A1(_2981_),
    .A2(_0405_),
    .B1(_0601_),
    .B2(_0409_),
    .Y(_1232_));
 sky130_fd_sc_hd__a221oi_1 _4518_ (.A1(_0981_),
    .A2(_3010_),
    .B1(_0982_),
    .B2(_0406_),
    .C1(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__nand2_1 _4519_ (.A(_0990_),
    .B(_0610_),
    .Y(_1234_));
 sky130_fd_sc_hd__nand2_1 _4520_ (.A(_0992_),
    .B(_3048_),
    .Y(_1235_));
 sky130_fd_sc_hd__nand2_1 _4521_ (.A(_1234_),
    .B(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__a221oi_1 _4522_ (.A1(_2943_),
    .A2(_0987_),
    .B1(_0841_),
    .B2(_0989_),
    .C1(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _4523_ (.A(_0428_),
    .B(_0657_),
    .Y(_1238_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_0999_),
    .B(_0926_),
    .Y(_1239_));
 sky130_fd_sc_hd__nand2_1 _4525_ (.A(_1238_),
    .B(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__a221oi_1 _4526_ (.A1(_0553_),
    .A2(_0996_),
    .B1(_2830_),
    .B2(_0997_),
    .C1(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__a22o_1 _4527_ (.A1(_0439_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[95] ),
    .B1(_0441_),
    .B2(_0638_),
    .X(_1242_));
 sky130_fd_sc_hd__o22ai_1 _4528_ (.A1(_3031_),
    .A2(_0446_),
    .B1(_0444_),
    .B2(_0449_),
    .Y(_1243_));
 sky130_fd_sc_hd__nor2_1 _4529_ (.A(_1242_),
    .B(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__and4_1 _4530_ (.A(_1233_),
    .B(_1237_),
    .C(_1241_),
    .D(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__and4_1 _4531_ (.A(_1206_),
    .B(_1222_),
    .C(_1231_),
    .D(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__nand3_1 _4532_ (.A(_1193_),
    .B(_0903_),
    .C(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__o21a_1 _4533_ (.A1(_2874_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1248_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_1247_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _4535_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(_1249_),
    .B(_1250_),
    .Y(_0299_));
 sky130_fd_sc_hd__a22o_1 _4537_ (.A1(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0777_),
    .X(_1251_));
 sky130_fd_sc_hd__a221oi_1 _4538_ (.A1(_1011_),
    .A2(_0781_),
    .B1(_3058_),
    .B2(_0782_),
    .C1(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_1 _4539_ (.A(_0791_),
    .B(_2990_),
    .Y(_1253_));
 sky130_fd_sc_hd__o21ai_1 _4540_ (.A1(_3154_),
    .A2(_0790_),
    .B1(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__a221oi_1 _4541_ (.A1(_3070_),
    .A2(_0787_),
    .B1(_2922_),
    .B2(_0788_),
    .C1(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__inv_2 _4542_ (.A(\egd_top.BitStream_buffer.BS_buffer[119] ),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _4543_ (.A(_0797_),
    .B(_2806_),
    .Y(_1257_));
 sky130_fd_sc_hd__o221a_1 _4544_ (.A1(_1256_),
    .A2(_3065_),
    .B1(_0538_),
    .B2(_0796_),
    .C1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__nand2_1 _4545_ (.A(_0802_),
    .B(_2800_),
    .Y(_1259_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(_0804_),
    .B(_2826_),
    .Y(_1260_));
 sky130_fd_sc_hd__nand2_1 _4547_ (.A(_1259_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__a221oi_1 _4548_ (.A1(_0330_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2818_),
    .C1(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__and4_1 _4549_ (.A(_1252_),
    .B(_1255_),
    .C(_1258_),
    .D(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__nand2_1 _4550_ (.A(_0812_),
    .B(_0402_),
    .Y(_1264_));
 sky130_fd_sc_hd__o21ai_1 _4551_ (.A1(_0859_),
    .A2(_0811_),
    .B1(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__a221oi_1 _4552_ (.A1(_2791_),
    .A2(_0810_),
    .B1(_3053_),
    .B2(_0809_),
    .C1(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_0818_),
    .B(_2822_),
    .Y(_1267_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(_0820_),
    .B(_2816_),
    .Y(_1268_));
 sky130_fd_sc_hd__nand2_1 _4555_ (.A(_1267_),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__a221oi_1 _4556_ (.A1(_0816_),
    .A2(_3066_),
    .B1(_0817_),
    .B2(_2824_),
    .C1(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__o22ai_1 _4557_ (.A1(_0984_),
    .A2(_0826_),
    .B1(_0601_),
    .B2(_0827_),
    .Y(_1271_));
 sky130_fd_sc_hd__a221oi_1 _4558_ (.A1(_0824_),
    .A2(_2913_),
    .B1(_0825_),
    .B2(_2980_),
    .C1(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__nand2_1 _4559_ (.A(_0833_),
    .B(_2814_),
    .Y(_1273_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_0835_),
    .B(_0458_),
    .Y(_1274_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_1273_),
    .B(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__a221oi_1 _4562_ (.A1(_0875_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2820_),
    .C1(_1275_),
    .Y(_1276_));
 sky130_fd_sc_hd__and4_1 _4563_ (.A(_1266_),
    .B(_1270_),
    .C(_1272_),
    .D(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_0844_),
    .B(_3034_),
    .Y(_1278_));
 sky130_fd_sc_hd__o21ai_1 _4565_ (.A1(_2944_),
    .A2(_0843_),
    .B1(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__a221oi_1 _4566_ (.A1(_0841_),
    .A2(_0840_),
    .B1(_2881_),
    .B2(_0842_),
    .C1(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__nand2_1 _4567_ (.A(_2867_),
    .B(_3090_),
    .Y(_1281_));
 sky130_fd_sc_hd__o21ai_1 _4568_ (.A1(_3078_),
    .A2(_0850_),
    .B1(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__a221oi_1 _4569_ (.A1(_2993_),
    .A2(_0848_),
    .B1(_3015_),
    .B2(_0849_),
    .C1(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__nand2_1 _4570_ (.A(_2858_),
    .B(_0495_),
    .Y(_1284_));
 sky130_fd_sc_hd__o21ai_1 _4571_ (.A1(_1005_),
    .A2(_2854_),
    .B1(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__a221oi_1 _4572_ (.A1(_0657_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_1000_),
    .C1(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__inv_2 _4573_ (.A(_0341_),
    .Y(_1287_));
 sky130_fd_sc_hd__o22ai_1 _4574_ (.A1(_1287_),
    .A2(_2912_),
    .B1(_0641_),
    .B2(_2917_),
    .Y(_1288_));
 sky130_fd_sc_hd__a221oi_1 _4575_ (.A1(_2907_),
    .A2(_0857_),
    .B1(_3127_),
    .B2(_0858_),
    .C1(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__and4_1 _4576_ (.A(_1280_),
    .B(_1283_),
    .C(_1286_),
    .D(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_0865_),
    .B(_3143_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2_1 _4578_ (.A(_0867_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _4579_ (.A(_1291_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__a221oi_1 _4580_ (.A1(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .A2(_0863_),
    .B1(_0864_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .C1(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__nand2_1 _4581_ (.A(_0874_),
    .B(_0583_),
    .Y(_1295_));
 sky130_fd_sc_hd__nand2_1 _4582_ (.A(_0877_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1296_));
 sky130_fd_sc_hd__nand2_1 _4583_ (.A(_1295_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__a221oi_1 _4584_ (.A1(_2904_),
    .A2(_0872_),
    .B1(_0830_),
    .B2(_0873_),
    .C1(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__nand2_1 _4585_ (.A(_0883_),
    .B(_1116_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _4586_ (.A(_0885_),
    .B(_0988_),
    .Y(_1300_));
 sky130_fd_sc_hd__inv_2 _4587_ (.A(\egd_top.BitStream_buffer.BS_buffer[67] ),
    .Y(_1301_));
 sky130_fd_sc_hd__or2_1 _4588_ (.A(_1301_),
    .B(_0889_),
    .X(_1302_));
 sky130_fd_sc_hd__o2111a_1 _4589_ (.A1(_3011_),
    .A2(_0882_),
    .B1(_1299_),
    .C1(_1300_),
    .D1(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__nand2_1 _4590_ (.A(_0895_),
    .B(_2828_),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(_0897_),
    .B(_0464_),
    .Y(_1305_));
 sky130_fd_sc_hd__nand2_1 _4592_ (.A(_1304_),
    .B(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__a221oi_1 _4593_ (.A1(_0892_),
    .A2(_2859_),
    .B1(_0893_),
    .B2(_0926_),
    .C1(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__and4_1 _4594_ (.A(_1294_),
    .B(_1298_),
    .C(_1303_),
    .D(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__and4_1 _4595_ (.A(_1263_),
    .B(_1277_),
    .C(_1290_),
    .D(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__o22ai_1 _4596_ (.A1(_0492_),
    .A2(_3131_),
    .B1(_0574_),
    .B2(_3135_),
    .Y(_1310_));
 sky130_fd_sc_hd__a221oi_1 _4597_ (.A1(_0343_),
    .A2(_3126_),
    .B1(_2974_),
    .B2(_3123_),
    .C1(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__nand2_1 _4598_ (.A(_3118_),
    .B(_3115_),
    .Y(_1312_));
 sky130_fd_sc_hd__o21ai_1 _4599_ (.A1(_2952_),
    .A2(_3110_),
    .B1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__a221oi_2 _4600_ (.A1(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .A2(_0907_),
    .B1(_3139_),
    .B2(_0908_),
    .C1(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__nand2_1 _4601_ (.A(_3100_),
    .B(_2887_),
    .Y(_1315_));
 sky130_fd_sc_hd__o21ai_1 _4602_ (.A1(_1171_),
    .A2(_3093_),
    .B1(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__a221oi_1 _4603_ (.A1(_2935_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_2848_),
    .C1(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__or2_1 _4604_ (.A(_3008_),
    .B(_3080_),
    .X(_1318_));
 sky130_fd_sc_hd__or2_1 _4605_ (.A(_0650_),
    .B(_3084_),
    .X(_1319_));
 sky130_fd_sc_hd__nand2_1 _4606_ (.A(_3087_),
    .B(_0389_),
    .Y(_1320_));
 sky130_fd_sc_hd__o2111a_1 _4607_ (.A1(_0904_),
    .A2(_3077_),
    .B1(_1318_),
    .C1(_1319_),
    .D1(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__and4_1 _4608_ (.A(_1311_),
    .B(_1314_),
    .C(_1317_),
    .D(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__or2b_1 _4609_ (.A(_0923_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[91] ),
    .X(_1323_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(_0925_),
    .B(_0587_),
    .Y(_1324_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_1323_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__a221oi_1 _4612_ (.A1(_0742_),
    .A2(_0921_),
    .B1(_0477_),
    .B2(_0922_),
    .C1(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__a22o_1 _4613_ (.A1(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_1327_));
 sky130_fd_sc_hd__a22o_1 _4614_ (.A1(_0933_),
    .A2(_0420_),
    .B1(_0934_),
    .B2(_0607_),
    .X(_1328_));
 sky130_fd_sc_hd__nor2_1 _4615_ (.A(_1327_),
    .B(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__nand2_1 _4616_ (.A(_0939_),
    .B(_0333_),
    .Y(_1330_));
 sky130_fd_sc_hd__nand2_1 _4617_ (.A(_0941_),
    .B(_3105_),
    .Y(_1331_));
 sky130_fd_sc_hd__nand2_1 _4618_ (.A(_1330_),
    .B(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__a221oi_1 _4619_ (.A1(_0937_),
    .A2(_0366_),
    .B1(_2957_),
    .B2(_0938_),
    .C1(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_0947_),
    .B(_3142_),
    .Y(_1334_));
 sky130_fd_sc_hd__nand2_1 _4621_ (.A(_0949_),
    .B(_0398_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_1 _4622_ (.A(_1334_),
    .B(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hd__a221oi_1 _4623_ (.A1(_2959_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_0336_),
    .C1(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__and4_1 _4624_ (.A(_1326_),
    .B(_1329_),
    .C(_1333_),
    .D(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__o22ai_1 _4625_ (.A1(_3031_),
    .A2(_0956_),
    .B1(_0698_),
    .B2(_0958_),
    .Y(_1339_));
 sky130_fd_sc_hd__a221oi_2 _4626_ (.A1(_2810_),
    .A2(_0954_),
    .B1(_2808_),
    .B2(_0955_),
    .C1(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__o22ai_1 _4627_ (.A1(_0731_),
    .A2(_0963_),
    .B1(_0347_),
    .B2(_0964_),
    .Y(_1341_));
 sky130_fd_sc_hd__a221oi_1 _4628_ (.A1(_0656_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_0371_),
    .C1(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__o22ai_1 _4629_ (.A1(_3129_),
    .A2(_0969_),
    .B1(_0730_),
    .B2(_0971_),
    .Y(_1343_));
 sky130_fd_sc_hd__a221oi_1 _4630_ (.A1(_0967_),
    .A2(_0886_),
    .B1(_0968_),
    .B2(_2874_),
    .C1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__o22ai_1 _4631_ (.A1(_0575_),
    .A2(_0976_),
    .B1(_0970_),
    .B2(_0977_),
    .Y(_1345_));
 sky130_fd_sc_hd__a221oi_1 _4632_ (.A1(_0974_),
    .A2(_3146_),
    .B1(_0975_),
    .B2(_3132_),
    .C1(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__and4_1 _4633_ (.A(_1340_),
    .B(_1342_),
    .C(_1344_),
    .D(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__o22ai_1 _4634_ (.A1(_0506_),
    .A2(_0405_),
    .B1(_0756_),
    .B2(_0409_),
    .Y(_1348_));
 sky130_fd_sc_hd__a221oi_1 _4635_ (.A1(_0981_),
    .A2(_0406_),
    .B1(_0982_),
    .B2(_3040_),
    .C1(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand2_1 _4636_ (.A(_0990_),
    .B(_0443_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _4637_ (.A(_0992_),
    .B(_3002_),
    .Y(_1351_));
 sky130_fd_sc_hd__nand2_1 _4638_ (.A(_1350_),
    .B(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__a221oi_1 _4639_ (.A1(_0412_),
    .A2(_0987_),
    .B1(_3101_),
    .B2(_0989_),
    .C1(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand2_1 _4640_ (.A(_0428_),
    .B(_0894_),
    .Y(_1354_));
 sky130_fd_sc_hd__nand2_1 _4641_ (.A(_0999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[86] ),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_1 _4642_ (.A(_1354_),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__a221oi_1 _4643_ (.A1(_0709_),
    .A2(_0996_),
    .B1(_0463_),
    .B2(_0997_),
    .C1(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__a22o_1 _4644_ (.A1(_0439_),
    .A2(_0638_),
    .B1(_0441_),
    .B2(_0610_),
    .X(_1358_));
 sky130_fd_sc_hd__o22ai_1 _4645_ (.A1(_0526_),
    .A2(_0446_),
    .B1(_0619_),
    .B2(_0449_),
    .Y(_1359_));
 sky130_fd_sc_hd__nor2_1 _4646_ (.A(_1358_),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__and4_1 _4647_ (.A(_1349_),
    .B(_1353_),
    .C(_1357_),
    .D(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__and4_1 _4648_ (.A(_1322_),
    .B(_1338_),
    .C(_1347_),
    .D(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__nand3_1 _4649_ (.A(_1309_),
    .B(_0903_),
    .C(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__o21a_1 _4650_ (.A1(_0469_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1364_));
 sky130_fd_sc_hd__nand2_1 _4651_ (.A(_1363_),
    .B(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__nand2_1 _4652_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_1366_));
 sky130_fd_sc_hd__nand2_1 _4653_ (.A(_1365_),
    .B(_1366_),
    .Y(_0298_));
 sky130_fd_sc_hd__a22o_1 _4654_ (.A1(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_1011_),
    .X(_1367_));
 sky130_fd_sc_hd__a221oi_1 _4655_ (.A1(_0886_),
    .A2(_0781_),
    .B1(_3066_),
    .B2(_0782_),
    .C1(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_0791_),
    .B(_3058_),
    .Y(_1369_));
 sky130_fd_sc_hd__o21ai_1 _4657_ (.A1(_0567_),
    .A2(_0790_),
    .B1(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__a221oi_1 _4658_ (.A1(_0330_),
    .A2(_0787_),
    .B1(_2913_),
    .B2(_0788_),
    .C1(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__inv_2 _4659_ (.A(\egd_top.BitStream_buffer.BS_buffer[120] ),
    .Y(_1372_));
 sky130_fd_sc_hd__nand2_1 _4660_ (.A(_0797_),
    .B(_2808_),
    .Y(_1373_));
 sky130_fd_sc_hd__o221a_1 _4661_ (.A1(_1372_),
    .A2(_3065_),
    .B1(_0698_),
    .B2(_0796_),
    .C1(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__nand2_1 _4662_ (.A(_0802_),
    .B(_2802_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_0804_),
    .B(_2828_),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_1 _4664_ (.A(_1375_),
    .B(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__a221oi_1 _4665_ (.A1(_2791_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2820_),
    .C1(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__and4_1 _4666_ (.A(_1368_),
    .B(_1371_),
    .C(_1374_),
    .D(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__nand2_1 _4667_ (.A(_0812_),
    .B(_2863_),
    .Y(_1380_));
 sky130_fd_sc_hd__o21ai_1 _4668_ (.A1(_1052_),
    .A2(_0811_),
    .B1(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__a221oi_1 _4669_ (.A1(_2800_),
    .A2(_0810_),
    .B1(_2990_),
    .B2(_0809_),
    .C1(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_0818_),
    .B(_2824_),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_1 _4671_ (.A(_0820_),
    .B(_2818_),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_1 _4672_ (.A(_1383_),
    .B(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__a221oi_1 _4673_ (.A1(_0816_),
    .A2(_3153_),
    .B1(_0817_),
    .B2(_2826_),
    .C1(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__o22ai_1 _4674_ (.A1(_0403_),
    .A2(_0826_),
    .B1(_0756_),
    .B2(_0827_),
    .Y(_1387_));
 sky130_fd_sc_hd__a221oi_1 _4675_ (.A1(_0824_),
    .A2(_2980_),
    .B1(_0825_),
    .B2(_3097_),
    .C1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__nand2_1 _4676_ (.A(_0833_),
    .B(_2816_),
    .Y(_1389_));
 sky130_fd_sc_hd__nand2_1 _4677_ (.A(_0835_),
    .B(_0625_),
    .Y(_1390_));
 sky130_fd_sc_hd__nand2_1 _4678_ (.A(_1389_),
    .B(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a221oi_1 _4679_ (.A1(_0587_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2822_),
    .C1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__and4_1 _4680_ (.A(_1382_),
    .B(_1386_),
    .C(_1388_),
    .D(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_0844_),
    .B(_3048_),
    .Y(_1394_));
 sky130_fd_sc_hd__o21ai_1 _4682_ (.A1(_0489_),
    .A2(_0843_),
    .B1(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__a221oi_1 _4683_ (.A1(_3101_),
    .A2(_0840_),
    .B1(_2943_),
    .B2(_0842_),
    .C1(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__nand2_1 _4684_ (.A(_2867_),
    .B(_2907_),
    .Y(_1397_));
 sky130_fd_sc_hd__o21ai_1 _4685_ (.A1(_0544_),
    .A2(_0850_),
    .B1(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__a221oi_2 _4686_ (.A1(_3010_),
    .A2(_0848_),
    .B1(_3017_),
    .B2(_0849_),
    .C1(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_2858_),
    .B(_0657_),
    .Y(_1400_));
 sky130_fd_sc_hd__o21ai_1 _4688_ (.A1(_1126_),
    .A2(_2854_),
    .B1(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__a221oi_1 _4689_ (.A1(_0894_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0830_),
    .C1(_1401_),
    .Y(_1402_));
 sky130_fd_sc_hd__inv_2 _4690_ (.A(\egd_top.BitStream_buffer.BS_buffer[39] ),
    .Y(_1403_));
 sky130_fd_sc_hd__o22ai_1 _4691_ (.A1(_1403_),
    .A2(_2912_),
    .B1(_0859_),
    .B2(_2917_),
    .Y(_1404_));
 sky130_fd_sc_hd__a221oi_1 _4692_ (.A1(_3127_),
    .A2(_0857_),
    .B1(_3124_),
    .B2(_0858_),
    .C1(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__and4_1 _4693_ (.A(_1396_),
    .B(_1399_),
    .C(_1402_),
    .D(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__nand2_1 _4694_ (.A(_0865_),
    .B(_0336_),
    .Y(_1407_));
 sky130_fd_sc_hd__nand2_1 _4695_ (.A(_0867_),
    .B(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .Y(_1408_));
 sky130_fd_sc_hd__nand2_1 _4696_ (.A(_1407_),
    .B(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__a221oi_2 _4697_ (.A1(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .A2(_0863_),
    .B1(_0864_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .C1(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hd__nand2_1 _4698_ (.A(_0874_),
    .B(_0871_),
    .Y(_1411_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(_0877_),
    .B(_2931_),
    .Y(_1412_));
 sky130_fd_sc_hd__nand2_1 _4700_ (.A(_1411_),
    .B(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__a221oi_1 _4701_ (.A1(_0477_),
    .A2(_0872_),
    .B1(_0926_),
    .B2(_0873_),
    .C1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand2_1 _4702_ (.A(_0883_),
    .B(_0841_),
    .Y(_1415_));
 sky130_fd_sc_hd__nand2_1 _4703_ (.A(_0885_),
    .B(_1116_),
    .Y(_1416_));
 sky130_fd_sc_hd__inv_2 _4704_ (.A(\egd_top.BitStream_buffer.BS_buffer[68] ),
    .Y(_1417_));
 sky130_fd_sc_hd__or2_1 _4705_ (.A(_1417_),
    .B(_0889_),
    .X(_1418_));
 sky130_fd_sc_hd__o2111a_1 _4706_ (.A1(_0407_),
    .A2(_0882_),
    .B1(_1415_),
    .C1(_1416_),
    .D1(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_0895_),
    .B(\egd_top.BitStream_buffer.BS_buffer[0] ),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _4708_ (.A(_0897_),
    .B(_2959_),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _4709_ (.A(_1420_),
    .B(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__a221oi_1 _4710_ (.A1(_0892_),
    .A2(_2830_),
    .B1(_0893_),
    .B2(_0920_),
    .C1(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__and4_1 _4711_ (.A(_1410_),
    .B(_1414_),
    .C(_1419_),
    .D(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__and4_1 _4712_ (.A(_1379_),
    .B(_1393_),
    .C(_1406_),
    .D(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__o22ai_1 _4713_ (.A1(_0653_),
    .A2(_3131_),
    .B1(_0730_),
    .B2(_3135_),
    .Y(_1426_));
 sky130_fd_sc_hd__a221oi_1 _4714_ (.A1(_2974_),
    .A2(_3126_),
    .B1(_0333_),
    .B2(_3123_),
    .C1(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_1 _4715_ (.A(_3118_),
    .B(_0385_),
    .Y(_1428_));
 sky130_fd_sc_hd__o21ai_1 _4716_ (.A1(_0492_),
    .A2(_3110_),
    .B1(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hd__a221oi_1 _4717_ (.A1(_3115_),
    .A2(_0907_),
    .B1(_0398_),
    .B2(_0908_),
    .C1(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_1 _4718_ (.A(_3100_),
    .B(_3007_),
    .Y(_1431_));
 sky130_fd_sc_hd__o21ai_1 _4719_ (.A1(_1287_),
    .A2(_3093_),
    .B1(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__a221oi_1 _4720_ (.A1(_0378_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_0464_),
    .C1(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__or2_1 _4721_ (.A(_0516_),
    .B(_3080_),
    .X(_1434_));
 sky130_fd_sc_hd__or2_1 _4722_ (.A(_0881_),
    .B(_3084_),
    .X(_1435_));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(_3087_),
    .B(_2951_),
    .Y(_1436_));
 sky130_fd_sc_hd__o2111a_1 _4724_ (.A1(_1075_),
    .A2(_3077_),
    .B1(_1434_),
    .C1(_1435_),
    .D1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__and4_1 _4725_ (.A(_1427_),
    .B(_1430_),
    .C(_1433_),
    .D(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__or2b_1 _4726_ (.A(_0923_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .X(_1439_));
 sky130_fd_sc_hd__nand2_1 _4727_ (.A(_0925_),
    .B(_0742_),
    .Y(_1440_));
 sky130_fd_sc_hd__nand2_1 _4728_ (.A(_1439_),
    .B(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__a221oi_1 _4729_ (.A1(_0638_),
    .A2(_0922_),
    .B1(_0583_),
    .B2(_0921_),
    .C1(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__a22o_1 _4730_ (.A1(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .X(_1443_));
 sky130_fd_sc_hd__a22o_1 _4731_ (.A1(_0933_),
    .A2(_0607_),
    .B1(_0934_),
    .B2(_2904_),
    .X(_1444_));
 sky130_fd_sc_hd__nor2_1 _4732_ (.A(_1443_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_0939_),
    .B(_3143_),
    .Y(_1446_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(_0941_),
    .B(_0553_),
    .Y(_1447_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_1446_),
    .B(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__a221oi_1 _4736_ (.A1(_0937_),
    .A2(_0435_),
    .B1(_0371_),
    .B2(_0938_),
    .C1(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__nand2_1 _4737_ (.A(_0947_),
    .B(_3139_),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0949_),
    .B(_0366_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(_1450_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__a221oi_1 _4740_ (.A1(_0495_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_3146_),
    .C1(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__and4_1 _4741_ (.A(_1442_),
    .B(_1445_),
    .C(_1449_),
    .D(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__o22ai_1 _4742_ (.A1(_0526_),
    .A2(_0956_),
    .B1(_0795_),
    .B2(_0958_),
    .Y(_1455_));
 sky130_fd_sc_hd__a221oi_2 _4743_ (.A1(_2812_),
    .A2(_0954_),
    .B1(_2810_),
    .B2(_0955_),
    .C1(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__o22ai_1 _4744_ (.A1(_0970_),
    .A2(_0963_),
    .B1(_0574_),
    .B2(_0964_),
    .Y(_1457_));
 sky130_fd_sc_hd__a221oi_1 _4745_ (.A1(_3105_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_0656_),
    .C1(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__o22ai_1 _4746_ (.A1(_0561_),
    .A2(_0969_),
    .B1(_3075_),
    .B2(_0971_),
    .Y(_1459_));
 sky130_fd_sc_hd__a221oi_1 _4747_ (.A1(_0967_),
    .A2(_2874_),
    .B1(_0968_),
    .B2(_0469_),
    .C1(_1459_),
    .Y(_1460_));
 sky130_fd_sc_hd__o22ai_1 _4748_ (.A1(_0731_),
    .A2(_0976_),
    .B1(_0347_),
    .B2(_0977_),
    .Y(_1461_));
 sky130_fd_sc_hd__a221oi_1 _4749_ (.A1(_0974_),
    .A2(_3132_),
    .B1(_0975_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .C1(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__and4_1 _4750_ (.A(_1456_),
    .B(_1458_),
    .C(_1460_),
    .D(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__o22ai_1 _4751_ (.A1(_3091_),
    .A2(_0405_),
    .B1(_0983_),
    .B2(_0409_),
    .Y(_1464_));
 sky130_fd_sc_hd__a221oi_1 _4752_ (.A1(_0981_),
    .A2(_3040_),
    .B1(_0982_),
    .B2(_3015_),
    .C1(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(_0990_),
    .B(_2987_),
    .Y(_1466_));
 sky130_fd_sc_hd__nand2_1 _4754_ (.A(_0992_),
    .B(_3030_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _4755_ (.A(_1466_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__a221oi_4 _4756_ (.A1(_0414_),
    .A2(_0987_),
    .B1(_0551_),
    .B2(_0989_),
    .C1(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_0428_),
    .B(_1000_),
    .Y(_1470_));
 sky130_fd_sc_hd__nand2_1 _4758_ (.A(_0999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[87] ),
    .Y(_1471_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(_1470_),
    .B(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__a221oi_1 _4760_ (.A1(_2859_),
    .A2(_0996_),
    .B1(_2848_),
    .B2(_0997_),
    .C1(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__a22o_1 _4761_ (.A1(_0439_),
    .A2(_0610_),
    .B1(_0441_),
    .B2(_0443_),
    .X(_1474_));
 sky130_fd_sc_hd__o22ai_1 _4762_ (.A1(_0686_),
    .A2(_0446_),
    .B1(_0772_),
    .B2(_0449_),
    .Y(_1475_));
 sky130_fd_sc_hd__nor2_1 _4763_ (.A(_1474_),
    .B(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__and4_1 _4764_ (.A(_1465_),
    .B(_1469_),
    .C(_1473_),
    .D(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__and4_1 _4765_ (.A(_1438_),
    .B(_1454_),
    .C(_1463_),
    .D(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__nand3_1 _4766_ (.A(_1425_),
    .B(_0903_),
    .C(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__o21a_1 _4767_ (.A1(_0988_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1480_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_1479_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__nand2_1 _4769_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2_1 _4770_ (.A(_1481_),
    .B(_1482_),
    .Y(_0297_));
 sky130_fd_sc_hd__a22o_1 _4771_ (.A1(\egd_top.BitStream_buffer.BS_buffer[3] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0886_),
    .X(_1483_));
 sky130_fd_sc_hd__a221oi_1 _4772_ (.A1(_2874_),
    .A2(_0781_),
    .B1(_3153_),
    .B2(_0782_),
    .C1(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__nand2_1 _4773_ (.A(_0791_),
    .B(_3066_),
    .Y(_1485_));
 sky130_fd_sc_hd__o21ai_1 _4774_ (.A1(_0723_),
    .A2(_0790_),
    .B1(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__a221oi_1 _4775_ (.A1(_2791_),
    .A2(_0787_),
    .B1(_2980_),
    .B2(_0788_),
    .C1(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__inv_2 _4776_ (.A(\egd_top.BitStream_buffer.BS_buffer[121] ),
    .Y(_1488_));
 sky130_fd_sc_hd__nand2_1 _4777_ (.A(_0797_),
    .B(_2810_),
    .Y(_1489_));
 sky130_fd_sc_hd__o221a_1 _4778_ (.A1(_1488_),
    .A2(_3065_),
    .B1(_0795_),
    .B2(_0796_),
    .C1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(_0802_),
    .B(_2804_),
    .Y(_1491_));
 sky130_fd_sc_hd__nand2_1 _4780_ (.A(_0804_),
    .B(_0458_),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_1491_),
    .B(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__a221oi_1 _4782_ (.A1(_2800_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2822_),
    .C1(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__and4_1 _4783_ (.A(_1484_),
    .B(_1487_),
    .C(_1490_),
    .D(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__nand2_1 _4784_ (.A(_0812_),
    .B(_2920_),
    .Y(_1496_));
 sky130_fd_sc_hd__o21ai_1 _4785_ (.A1(_1171_),
    .A2(_0811_),
    .B1(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__a221oi_1 _4786_ (.A1(_2802_),
    .A2(_0810_),
    .B1(_3058_),
    .B2(_0809_),
    .C1(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2_1 _4787_ (.A(_0818_),
    .B(_2826_),
    .Y(_1499_));
 sky130_fd_sc_hd__nand2_1 _4788_ (.A(_0820_),
    .B(_2820_),
    .Y(_1500_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_1499_),
    .B(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__a221oi_1 _4790_ (.A1(_0816_),
    .A2(_3070_),
    .B1(_0817_),
    .B2(_2828_),
    .C1(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__o22ai_1 _4791_ (.A1(_0601_),
    .A2(_0826_),
    .B1(_0983_),
    .B2(_0827_),
    .Y(_1503_));
 sky130_fd_sc_hd__a221oi_1 _4792_ (.A1(_0824_),
    .A2(_3097_),
    .B1(_0825_),
    .B2(_3090_),
    .C1(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_0833_),
    .B(_2818_),
    .Y(_1505_));
 sky130_fd_sc_hd__nand2_1 _4794_ (.A(_0835_),
    .B(_0777_),
    .Y(_1506_));
 sky130_fd_sc_hd__nand2_1 _4795_ (.A(_1505_),
    .B(_1506_),
    .Y(_1507_));
 sky130_fd_sc_hd__a221oi_2 _4796_ (.A1(_0742_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2824_),
    .C1(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__and4_1 _4797_ (.A(_1498_),
    .B(_1502_),
    .C(_1504_),
    .D(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__nand2_1 _4798_ (.A(_0844_),
    .B(_3002_),
    .Y(_1510_));
 sky130_fd_sc_hd__o21ai_1 _4799_ (.A1(_0650_),
    .A2(_0843_),
    .B1(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__a221oi_1 _4800_ (.A1(_0551_),
    .A2(_0840_),
    .B1(_0412_),
    .B2(_0842_),
    .C1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand2_1 _4801_ (.A(_2867_),
    .B(_3127_),
    .Y(_1513_));
 sky130_fd_sc_hd__o21ai_1 _4802_ (.A1(_2944_),
    .A2(_0850_),
    .B1(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__a221oi_1 _4803_ (.A1(_0406_),
    .A2(_0848_),
    .B1(_0402_),
    .B2(_0849_),
    .C1(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__nand2_1 _4804_ (.A(_2858_),
    .B(_0894_),
    .Y(_1516_));
 sky130_fd_sc_hd__o21ai_1 _4805_ (.A1(_3031_),
    .A2(_2854_),
    .B1(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__a221oi_1 _4806_ (.A1(_1000_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0926_),
    .C1(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__inv_2 _4807_ (.A(\egd_top.BitStream_buffer.BS_buffer[40] ),
    .Y(_1519_));
 sky130_fd_sc_hd__o22ai_1 _4808_ (.A1(_1519_),
    .A2(_2912_),
    .B1(_1052_),
    .B2(_2917_),
    .Y(_1520_));
 sky130_fd_sc_hd__a221oi_1 _4809_ (.A1(_3124_),
    .A2(_0857_),
    .B1(_0395_),
    .B2(_0858_),
    .C1(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__and4_1 _4810_ (.A(_1512_),
    .B(_1515_),
    .C(_1518_),
    .D(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__nand2_1 _4811_ (.A(_0865_),
    .B(_3146_),
    .Y(_1523_));
 sky130_fd_sc_hd__nand2_1 _4812_ (.A(_0867_),
    .B(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .Y(_1524_));
 sky130_fd_sc_hd__nand2_1 _4813_ (.A(_1523_),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__a221oi_2 _4814_ (.A1(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .A2(_0863_),
    .B1(_0864_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .C1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _4815_ (.A(_0874_),
    .B(_0420_),
    .Y(_1527_));
 sky130_fd_sc_hd__nand2_1 _4816_ (.A(_0877_),
    .B(_2939_),
    .Y(_1528_));
 sky130_fd_sc_hd__nand2_1 _4817_ (.A(_1527_),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__a221oi_1 _4818_ (.A1(_0638_),
    .A2(_0872_),
    .B1(_0920_),
    .B2(_0873_),
    .C1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__nand2_1 _4819_ (.A(_0883_),
    .B(_3101_),
    .Y(_1531_));
 sky130_fd_sc_hd__nand2_1 _4820_ (.A(_0885_),
    .B(_0841_),
    .Y(_1532_));
 sky130_fd_sc_hd__inv_2 _4821_ (.A(\egd_top.BitStream_buffer.BS_buffer[69] ),
    .Y(_1533_));
 sky130_fd_sc_hd__or2_1 _4822_ (.A(_1533_),
    .B(_0889_),
    .X(_1534_));
 sky130_fd_sc_hd__o2111a_1 _4823_ (.A1(_0602_),
    .A2(_0882_),
    .B1(_1531_),
    .C1(_1532_),
    .D1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__nand2_1 _4824_ (.A(_0895_),
    .B(\egd_top.BitStream_buffer.BS_buffer[1] ),
    .Y(_1536_));
 sky130_fd_sc_hd__nand2_1 _4825_ (.A(_0897_),
    .B(_0495_),
    .Y(_1537_));
 sky130_fd_sc_hd__nand2_1 _4826_ (.A(_1536_),
    .B(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__a221oi_1 _4827_ (.A1(_0892_),
    .A2(_0463_),
    .B1(_0893_),
    .B2(_0875_),
    .C1(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__and4_1 _4828_ (.A(_1526_),
    .B(_1530_),
    .C(_1535_),
    .D(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__and4_1 _4829_ (.A(_1495_),
    .B(_1509_),
    .C(_1522_),
    .D(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__o22ai_1 _4830_ (.A1(_0888_),
    .A2(_3131_),
    .B1(_3075_),
    .B2(_3135_),
    .Y(_1542_));
 sky130_fd_sc_hd__a221oi_1 _4831_ (.A1(_0333_),
    .A2(_3126_),
    .B1(_3143_),
    .B2(_3123_),
    .C1(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_3118_),
    .B(_0389_),
    .Y(_1544_));
 sky130_fd_sc_hd__o21ai_1 _4833_ (.A1(_0653_),
    .A2(_3110_),
    .B1(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__a221oi_1 _4834_ (.A1(_0385_),
    .A2(_0907_),
    .B1(_0366_),
    .B2(_0908_),
    .C1(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__nand2_1 _4835_ (.A(_3100_),
    .B(_2993_),
    .Y(_1547_));
 sky130_fd_sc_hd__o21ai_1 _4836_ (.A1(_1403_),
    .A2(_3093_),
    .B1(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__a221oi_2 _4837_ (.A1(_0341_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_2959_),
    .C1(_1548_),
    .Y(_1549_));
 sky130_fd_sc_hd__or2_1 _4838_ (.A(_3011_),
    .B(_3080_),
    .X(_1550_));
 sky130_fd_sc_hd__or2_1 _4839_ (.A(_3008_),
    .B(_3084_),
    .X(_1551_));
 sky130_fd_sc_hd__nand2_1 _4840_ (.A(_3087_),
    .B(_0392_),
    .Y(_1552_));
 sky130_fd_sc_hd__o2111a_1 _4841_ (.A1(_2952_),
    .A2(_3077_),
    .B1(_1550_),
    .C1(_1551_),
    .D1(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__and4_1 _4842_ (.A(_1543_),
    .B(_1546_),
    .C(_1549_),
    .D(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__o22ai_1 _4843_ (.A1(_0686_),
    .A2(_0956_),
    .B1(_1021_),
    .B2(_0958_),
    .Y(_1555_));
 sky130_fd_sc_hd__a221oi_2 _4844_ (.A1(_2814_),
    .A2(_0954_),
    .B1(_2812_),
    .B2(_0955_),
    .C1(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__o22ai_1 _4845_ (.A1(_0347_),
    .A2(_0963_),
    .B1(_0730_),
    .B2(_0964_),
    .Y(_1557_));
 sky130_fd_sc_hd__a221oi_1 _4846_ (.A1(_0553_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_3105_),
    .C1(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__o22ai_1 _4847_ (.A1(_0717_),
    .A2(_0969_),
    .B1(_0543_),
    .B2(_0971_),
    .Y(_1559_));
 sky130_fd_sc_hd__a221oi_1 _4848_ (.A1(_0967_),
    .A2(_0469_),
    .B1(_0968_),
    .B2(_0988_),
    .C1(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__o22ai_1 _4849_ (.A1(_0970_),
    .A2(_0976_),
    .B1(_0574_),
    .B2(_0977_),
    .Y(_1561_));
 sky130_fd_sc_hd__a221oi_1 _4850_ (.A1(_0974_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .B1(_0975_),
    .B2(_2931_),
    .C1(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__and4_1 _4851_ (.A(_1556_),
    .B(_1558_),
    .C(_1560_),
    .D(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__o22ai_1 _4852_ (.A1(_2908_),
    .A2(_0405_),
    .B1(_2914_),
    .B2(_0409_),
    .Y(_1564_));
 sky130_fd_sc_hd__a221oi_1 _4853_ (.A1(_0981_),
    .A2(_3015_),
    .B1(_0982_),
    .B2(_3017_),
    .C1(_1564_),
    .Y(_1565_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_0990_),
    .B(_3034_),
    .Y(_1566_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_0992_),
    .B(_3037_),
    .Y(_1567_));
 sky130_fd_sc_hd__nand2_1 _4856_ (.A(_1566_),
    .B(_1567_),
    .Y(_1568_));
 sky130_fd_sc_hd__a221oi_1 _4857_ (.A1(_2887_),
    .A2(_0987_),
    .B1(_2881_),
    .B2(_0989_),
    .C1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hd__nand2_1 _4858_ (.A(_0428_),
    .B(_0830_),
    .Y(_1570_));
 sky130_fd_sc_hd__nand2_1 _4859_ (.A(_0999_),
    .B(_0587_),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_1 _4860_ (.A(_1570_),
    .B(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__a221oi_1 _4861_ (.A1(_2830_),
    .A2(_0996_),
    .B1(_0464_),
    .B2(_0997_),
    .C1(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hd__a22o_1 _4862_ (.A1(_0439_),
    .A2(_0443_),
    .B1(_0441_),
    .B2(_2987_),
    .X(_1574_));
 sky130_fd_sc_hd__o22ai_1 _4863_ (.A1(_0789_),
    .A2(_0446_),
    .B1(_1005_),
    .B2(_0449_),
    .Y(_1575_));
 sky130_fd_sc_hd__nor2_1 _4864_ (.A(_1574_),
    .B(_1575_),
    .Y(_1576_));
 sky130_fd_sc_hd__and4_1 _4865_ (.A(_1565_),
    .B(_1569_),
    .C(_1573_),
    .D(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__nand2_1 _4866_ (.A(_0925_),
    .B(_0583_),
    .Y(_1578_));
 sky130_fd_sc_hd__o21ai_1 _4867_ (.A1(_0447_),
    .A2(_0923_),
    .B1(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__a221oi_1 _4868_ (.A1(_0610_),
    .A2(_0922_),
    .B1(_0871_),
    .B2(_0921_),
    .C1(_1579_),
    .Y(_1580_));
 sky130_fd_sc_hd__nand2_1 _4869_ (.A(_0947_),
    .B(_0398_),
    .Y(_1581_));
 sky130_fd_sc_hd__nand2_1 _4870_ (.A(_0949_),
    .B(_0435_),
    .Y(_1582_));
 sky130_fd_sc_hd__nand2_1 _4871_ (.A(_1581_),
    .B(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__a221oi_1 _4872_ (.A1(_0657_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_3132_),
    .C1(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__nand2_1 _4873_ (.A(_0939_),
    .B(_0336_),
    .Y(_1585_));
 sky130_fd_sc_hd__nand2_1 _4874_ (.A(_0941_),
    .B(_0709_),
    .Y(_1586_));
 sky130_fd_sc_hd__nand2_1 _4875_ (.A(_1585_),
    .B(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__a221oi_2 _4876_ (.A1(_0937_),
    .A2(_2957_),
    .B1(_0656_),
    .B2(_0938_),
    .C1(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__a22o_1 _4877_ (.A1(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .X(_1589_));
 sky130_fd_sc_hd__a22o_1 _4878_ (.A1(_0933_),
    .A2(_2904_),
    .B1(_0934_),
    .B2(_0477_),
    .X(_1590_));
 sky130_fd_sc_hd__nor2_1 _4879_ (.A(_1589_),
    .B(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__and4_1 _4880_ (.A(_1580_),
    .B(_1584_),
    .C(_1588_),
    .D(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__and4_1 _4881_ (.A(_1554_),
    .B(_1563_),
    .C(_1577_),
    .D(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__nand3_1 _4882_ (.A(_1541_),
    .B(_0903_),
    .C(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__o21a_1 _4883_ (.A1(_1116_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1595_));
 sky130_fd_sc_hd__nand2_1 _4884_ (.A(_1594_),
    .B(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_1 _4886_ (.A(_1596_),
    .B(_1597_),
    .Y(_0296_));
 sky130_fd_sc_hd__a22o_1 _4887_ (.A1(\egd_top.BitStream_buffer.BS_buffer[4] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_2874_),
    .X(_1598_));
 sky130_fd_sc_hd__a221oi_2 _4888_ (.A1(_0469_),
    .A2(_0781_),
    .B1(_3070_),
    .B2(_0782_),
    .C1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__nand2_1 _4889_ (.A(_0791_),
    .B(_3153_),
    .Y(_1600_));
 sky130_fd_sc_hd__o21ai_1 _4890_ (.A1(_0957_),
    .A2(_0790_),
    .B1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__a221oi_1 _4891_ (.A1(_2800_),
    .A2(_0787_),
    .B1(_3097_),
    .B2(_0788_),
    .C1(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__inv_2 _4892_ (.A(\egd_top.BitStream_buffer.BS_buffer[122] ),
    .Y(_1603_));
 sky130_fd_sc_hd__nand2_1 _4893_ (.A(_0797_),
    .B(_2812_),
    .Y(_1604_));
 sky130_fd_sc_hd__o221a_1 _4894_ (.A1(_1603_),
    .A2(_3065_),
    .B1(_1021_),
    .B2(_0796_),
    .C1(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__nand2_1 _4895_ (.A(_0802_),
    .B(_2806_),
    .Y(_1606_));
 sky130_fd_sc_hd__nand2_1 _4896_ (.A(_0804_),
    .B(_0625_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand2_1 _4897_ (.A(_1606_),
    .B(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__a221oi_1 _4898_ (.A1(_2802_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2824_),
    .C1(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__and4_1 _4899_ (.A(_1599_),
    .B(_1602_),
    .C(_1605_),
    .D(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__nand2_1 _4900_ (.A(_0812_),
    .B(_2922_),
    .Y(_1611_));
 sky130_fd_sc_hd__o21ai_1 _4901_ (.A1(_1287_),
    .A2(_0811_),
    .B1(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__a221oi_1 _4902_ (.A1(_2804_),
    .A2(_0810_),
    .B1(_3066_),
    .B2(_0809_),
    .C1(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__nand2_1 _4903_ (.A(_0818_),
    .B(_2828_),
    .Y(_1614_));
 sky130_fd_sc_hd__nand2_1 _4904_ (.A(_0820_),
    .B(_2822_),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_1614_),
    .B(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__a221oi_1 _4906_ (.A1(_0816_),
    .A2(_0330_),
    .B1(_0817_),
    .B2(_0458_),
    .C1(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__o22ai_1 _4907_ (.A1(_0756_),
    .A2(_0826_),
    .B1(_2914_),
    .B2(_0827_),
    .Y(_1618_));
 sky130_fd_sc_hd__a221oi_1 _4908_ (.A1(_0824_),
    .A2(_3090_),
    .B1(_0825_),
    .B2(_2907_),
    .C1(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__nand2_1 _4909_ (.A(_0833_),
    .B(_2820_),
    .Y(_1620_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(_0835_),
    .B(_1011_),
    .Y(_1621_));
 sky130_fd_sc_hd__nand2_1 _4911_ (.A(_1620_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__a221oi_1 _4912_ (.A1(_0583_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2826_),
    .C1(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__and4_1 _4913_ (.A(_1613_),
    .B(_1617_),
    .C(_1619_),
    .D(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_1 _4914_ (.A(_0844_),
    .B(_3030_),
    .Y(_1625_));
 sky130_fd_sc_hd__o21ai_1 _4915_ (.A1(_0881_),
    .A2(_0843_),
    .B1(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__a221oi_1 _4916_ (.A1(_2881_),
    .A2(_0840_),
    .B1(_0414_),
    .B2(_0842_),
    .C1(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__nand2_1 _4917_ (.A(_2867_),
    .B(_3124_),
    .Y(_1628_));
 sky130_fd_sc_hd__o21ai_1 _4918_ (.A1(_0489_),
    .A2(_0850_),
    .B1(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__a221oi_1 _4919_ (.A1(_3040_),
    .A2(_0848_),
    .B1(_2863_),
    .B2(_0849_),
    .C1(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__nand2_1 _4920_ (.A(_2858_),
    .B(_1000_),
    .Y(_1631_));
 sky130_fd_sc_hd__o21ai_1 _4921_ (.A1(_0526_),
    .A2(_2854_),
    .B1(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__a221oi_1 _4922_ (.A1(_0830_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0920_),
    .C1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__o22ai_1 _4923_ (.A1(_0334_),
    .A2(_2912_),
    .B1(_1171_),
    .B2(_2917_),
    .Y(_1634_));
 sky130_fd_sc_hd__a221oi_1 _4924_ (.A1(_0395_),
    .A2(_0857_),
    .B1(_2935_),
    .B2(_0858_),
    .C1(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__and4_1 _4925_ (.A(_1627_),
    .B(_1630_),
    .C(_1633_),
    .D(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__nand2_1 _4926_ (.A(_0865_),
    .B(_3132_),
    .Y(_1637_));
 sky130_fd_sc_hd__nand2_1 _4927_ (.A(_0867_),
    .B(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .Y(_1638_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_1637_),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__a221oi_2 _4929_ (.A1(_3115_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .C1(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_0874_),
    .B(_0607_),
    .Y(_1641_));
 sky130_fd_sc_hd__nand2_1 _4931_ (.A(_0877_),
    .B(_2926_),
    .Y(_1642_));
 sky130_fd_sc_hd__nand2_1 _4932_ (.A(_1641_),
    .B(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__a221oi_1 _4933_ (.A1(_0610_),
    .A2(_0872_),
    .B1(_0875_),
    .B2(_0873_),
    .C1(_1643_),
    .Y(_1644_));
 sky130_fd_sc_hd__nand2_1 _4934_ (.A(_0883_),
    .B(_0551_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand2_1 _4935_ (.A(_0885_),
    .B(_3101_),
    .Y(_1646_));
 sky130_fd_sc_hd__inv_2 _4936_ (.A(\egd_top.BitStream_buffer.BS_buffer[70] ),
    .Y(_1647_));
 sky130_fd_sc_hd__or2_1 _4937_ (.A(_1647_),
    .B(_0889_),
    .X(_1648_));
 sky130_fd_sc_hd__o2111a_1 _4938_ (.A1(_0757_),
    .A2(_0882_),
    .B1(_1645_),
    .C1(_1646_),
    .D1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__nand2_1 _4939_ (.A(_0895_),
    .B(\egd_top.BitStream_buffer.BS_buffer[2] ),
    .Y(_1650_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(_0897_),
    .B(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .Y(_1651_));
 sky130_fd_sc_hd__nand2_1 _4941_ (.A(_1650_),
    .B(_1651_),
    .Y(_1652_));
 sky130_fd_sc_hd__a221oi_1 _4942_ (.A1(_0892_),
    .A2(_2848_),
    .B1(_0893_),
    .B2(_0587_),
    .C1(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__and4_1 _4943_ (.A(_1640_),
    .B(_1644_),
    .C(_1649_),
    .D(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__and4_1 _4944_ (.A(_1610_),
    .B(_1624_),
    .C(_1636_),
    .D(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__o22ai_1 _4945_ (.A1(_1066_),
    .A2(_3131_),
    .B1(_0543_),
    .B2(_3135_),
    .Y(_1656_));
 sky130_fd_sc_hd__a221oi_1 _4946_ (.A1(_3143_),
    .A2(_3126_),
    .B1(_0336_),
    .B2(_3123_),
    .C1(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__nand2_1 _4947_ (.A(_3118_),
    .B(_2951_),
    .Y(_1658_));
 sky130_fd_sc_hd__o21ai_1 _4948_ (.A1(_0888_),
    .A2(_3110_),
    .B1(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__a221oi_2 _4949_ (.A1(_0389_),
    .A2(_0907_),
    .B1(_0435_),
    .B2(_0908_),
    .C1(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand2_1 _4950_ (.A(_3100_),
    .B(_3010_),
    .Y(_1661_));
 sky130_fd_sc_hd__o21ai_1 _4951_ (.A1(_1519_),
    .A2(_3093_),
    .B1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__a221oi_2 _4952_ (.A1(_0343_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_0495_),
    .C1(_1662_),
    .Y(_1663_));
 sky130_fd_sc_hd__or2_1 _4953_ (.A(_0407_),
    .B(_3080_),
    .X(_1664_));
 sky130_fd_sc_hd__or2_1 _4954_ (.A(_0516_),
    .B(_3084_),
    .X(_1665_));
 sky130_fd_sc_hd__nand2_1 _4955_ (.A(_3087_),
    .B(_3142_),
    .Y(_1666_));
 sky130_fd_sc_hd__o2111a_1 _4956_ (.A1(_0492_),
    .A2(_3077_),
    .B1(_1664_),
    .C1(_1665_),
    .D1(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__and4_1 _4957_ (.A(_1657_),
    .B(_1660_),
    .C(_1663_),
    .D(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__o22ai_2 _4958_ (.A1(_0789_),
    .A2(_0956_),
    .B1(_1140_),
    .B2(_0958_),
    .Y(_1669_));
 sky130_fd_sc_hd__a221oi_4 _4959_ (.A1(_2816_),
    .A2(_0954_),
    .B1(_2814_),
    .B2(_0955_),
    .C1(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__o22ai_1 _4960_ (.A1(_0574_),
    .A2(_0963_),
    .B1(_3075_),
    .B2(_0964_),
    .Y(_1671_));
 sky130_fd_sc_hd__a221oi_1 _4961_ (.A1(_0709_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_0553_),
    .C1(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__o22ai_1 _4962_ (.A1(_0904_),
    .A2(_0969_),
    .B1(_3108_),
    .B2(_0971_),
    .Y(_1673_));
 sky130_fd_sc_hd__a221oi_1 _4963_ (.A1(_0967_),
    .A2(_0988_),
    .B1(_0968_),
    .B2(_1116_),
    .C1(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hd__o22ai_1 _4964_ (.A1(_0347_),
    .A2(_0976_),
    .B1(_0730_),
    .B2(_0977_),
    .Y(_1675_));
 sky130_fd_sc_hd__a221oi_1 _4965_ (.A1(_0974_),
    .A2(_2931_),
    .B1(_0975_),
    .B2(_2939_),
    .C1(_1675_),
    .Y(_1676_));
 sky130_fd_sc_hd__and4_1 _4966_ (.A(_1670_),
    .B(_1672_),
    .C(_1674_),
    .D(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__o22ai_1 _4967_ (.A1(_0480_),
    .A2(_0405_),
    .B1(_2981_),
    .B2(_0409_),
    .Y(_1678_));
 sky130_fd_sc_hd__a221oi_1 _4968_ (.A1(_0981_),
    .A2(_3017_),
    .B1(_0982_),
    .B2(_0402_),
    .C1(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_0990_),
    .B(_3048_),
    .Y(_1680_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_0992_),
    .B(_3053_),
    .Y(_1681_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_1680_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__a221oi_1 _4972_ (.A1(_3007_),
    .A2(_0987_),
    .B1(_2943_),
    .B2(_0989_),
    .C1(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__nand2_1 _4973_ (.A(_0428_),
    .B(_0926_),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_1 _4974_ (.A(_0999_),
    .B(_0742_),
    .Y(_1685_));
 sky130_fd_sc_hd__nand2_1 _4975_ (.A(_1684_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__a221oi_1 _4976_ (.A1(_0463_),
    .A2(_0996_),
    .B1(_2959_),
    .B2(_0997_),
    .C1(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__a22o_1 _4977_ (.A1(_0439_),
    .A2(_2987_),
    .B1(_0441_),
    .B2(_3034_),
    .X(_1688_));
 sky130_fd_sc_hd__o22ai_1 _4978_ (.A1(_1017_),
    .A2(_0446_),
    .B1(_1126_),
    .B2(_0449_),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_1 _4979_ (.A(_1688_),
    .B(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__and4_1 _4980_ (.A(_1679_),
    .B(_1683_),
    .C(_1687_),
    .D(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__nand2_1 _4981_ (.A(_0925_),
    .B(_0871_),
    .Y(_1692_));
 sky130_fd_sc_hd__o21ai_1 _4982_ (.A1(_0620_),
    .A2(_0923_),
    .B1(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__a221oi_1 _4983_ (.A1(_0443_),
    .A2(_0922_),
    .B1(_0420_),
    .B2(_0921_),
    .C1(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__nand2_1 _4984_ (.A(_0947_),
    .B(_0366_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand2_1 _4985_ (.A(_0949_),
    .B(_2957_),
    .Y(_1696_));
 sky130_fd_sc_hd__nand2_1 _4986_ (.A(_1695_),
    .B(_1696_),
    .Y(_1697_));
 sky130_fd_sc_hd__a221oi_1 _4987_ (.A1(_0894_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .C1(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_0939_),
    .B(_3146_),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_1 _4989_ (.A(_0941_),
    .B(_2859_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand2_1 _4990_ (.A(_1699_),
    .B(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__a221oi_1 _4991_ (.A1(_0937_),
    .A2(_0371_),
    .B1(_3105_),
    .B2(_0938_),
    .C1(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__a22o_1 _4992_ (.A1(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .X(_1703_));
 sky130_fd_sc_hd__a22o_1 _4993_ (.A1(_0933_),
    .A2(_0477_),
    .B1(_0934_),
    .B2(_0638_),
    .X(_1704_));
 sky130_fd_sc_hd__nor2_1 _4994_ (.A(_1703_),
    .B(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__and4_2 _4995_ (.A(_1694_),
    .B(_1698_),
    .C(_1702_),
    .D(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__and4_1 _4996_ (.A(_1668_),
    .B(_1677_),
    .C(_1691_),
    .D(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__nand3_1 _4997_ (.A(_1655_),
    .B(_0903_),
    .C(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__o21a_1 _4998_ (.A1(_0841_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1709_));
 sky130_fd_sc_hd__nand2_1 _4999_ (.A(_1708_),
    .B(_1709_),
    .Y(_1710_));
 sky130_fd_sc_hd__nand2_1 _5000_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_1711_));
 sky130_fd_sc_hd__nand2_1 _5001_ (.A(_1710_),
    .B(_1711_),
    .Y(_0295_));
 sky130_fd_sc_hd__a22o_1 _5002_ (.A1(\egd_top.BitStream_buffer.BS_buffer[5] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0469_),
    .X(_1712_));
 sky130_fd_sc_hd__a221oi_1 _5003_ (.A1(_0988_),
    .A2(_0781_),
    .B1(_0330_),
    .B2(_0782_),
    .C1(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__nand2_1 _5004_ (.A(_0791_),
    .B(_3070_),
    .Y(_1714_));
 sky130_fd_sc_hd__o21ai_1 _5005_ (.A1(_3064_),
    .A2(_0790_),
    .B1(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__a221oi_1 _5006_ (.A1(_2802_),
    .A2(_0787_),
    .B1(_3090_),
    .B2(_0788_),
    .C1(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__inv_2 _5007_ (.A(\egd_top.BitStream_buffer.BS_buffer[123] ),
    .Y(_1717_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_0797_),
    .B(_2814_),
    .Y(_1718_));
 sky130_fd_sc_hd__o221a_1 _5009_ (.A1(_1717_),
    .A2(_3065_),
    .B1(_1140_),
    .B2(_0796_),
    .C1(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(_0802_),
    .B(_2808_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand2_1 _5011_ (.A(_0804_),
    .B(_0777_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand2_1 _5012_ (.A(_1720_),
    .B(_1721_),
    .Y(_1722_));
 sky130_fd_sc_hd__a221oi_1 _5013_ (.A1(_2804_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2826_),
    .C1(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__and4_1 _5014_ (.A(_1713_),
    .B(_1716_),
    .C(_1719_),
    .D(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_1 _5015_ (.A(_0812_),
    .B(_2913_),
    .Y(_1725_));
 sky130_fd_sc_hd__o21ai_1 _5016_ (.A1(_1403_),
    .A2(_0811_),
    .B1(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__a221oi_1 _5017_ (.A1(_2806_),
    .A2(_0810_),
    .B1(_3153_),
    .B2(_0809_),
    .C1(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__nand2_1 _5018_ (.A(_0818_),
    .B(_0458_),
    .Y(_1728_));
 sky130_fd_sc_hd__nand2_1 _5019_ (.A(_0820_),
    .B(_2824_),
    .Y(_1729_));
 sky130_fd_sc_hd__nand2_1 _5020_ (.A(_1728_),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__a221oi_1 _5021_ (.A1(_0816_),
    .A2(_2791_),
    .B1(_0817_),
    .B2(_0625_),
    .C1(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__o22ai_1 _5022_ (.A1(_0983_),
    .A2(_0826_),
    .B1(_2981_),
    .B2(_0827_),
    .Y(_1732_));
 sky130_fd_sc_hd__a221oi_1 _5023_ (.A1(_0824_),
    .A2(_2907_),
    .B1(_0825_),
    .B2(_3127_),
    .C1(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(_0833_),
    .B(_2822_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _5025_ (.A(_0835_),
    .B(_0886_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_1 _5026_ (.A(_1734_),
    .B(_1735_),
    .Y(_1736_));
 sky130_fd_sc_hd__a221oi_1 _5027_ (.A1(_0871_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_2828_),
    .C1(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__and4_1 _5028_ (.A(_1727_),
    .B(_1731_),
    .C(_1733_),
    .D(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__nand2_1 _5029_ (.A(_0844_),
    .B(_3037_),
    .Y(_1739_));
 sky130_fd_sc_hd__o21ai_1 _5030_ (.A1(_3008_),
    .A2(_0843_),
    .B1(_1739_),
    .Y(_1740_));
 sky130_fd_sc_hd__a221oi_1 _5031_ (.A1(_2943_),
    .A2(_0840_),
    .B1(_2887_),
    .B2(_0842_),
    .C1(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hd__nand2_1 _5032_ (.A(_2867_),
    .B(_0395_),
    .Y(_1742_));
 sky130_fd_sc_hd__o21ai_1 _5033_ (.A1(_0650_),
    .A2(_0850_),
    .B1(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hd__a221oi_1 _5034_ (.A1(_3015_),
    .A2(_0848_),
    .B1(_2920_),
    .B2(_0849_),
    .C1(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_2858_),
    .B(_0830_),
    .Y(_1745_));
 sky130_fd_sc_hd__o21ai_1 _5036_ (.A1(_0686_),
    .A2(_2854_),
    .B1(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__a221oi_1 _5037_ (.A1(_0926_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0875_),
    .C1(_1746_),
    .Y(_1747_));
 sky130_fd_sc_hd__o22ai_1 _5038_ (.A1(_3144_),
    .A2(_2912_),
    .B1(_1287_),
    .B2(_2917_),
    .Y(_1748_));
 sky130_fd_sc_hd__a221oi_1 _5039_ (.A1(_2935_),
    .A2(_0857_),
    .B1(_0378_),
    .B2(_0858_),
    .C1(_1748_),
    .Y(_1749_));
 sky130_fd_sc_hd__and4_1 _5040_ (.A(_1741_),
    .B(_1744_),
    .C(_1747_),
    .D(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__nand2_1 _5041_ (.A(_0865_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1751_));
 sky130_fd_sc_hd__nand2_1 _5042_ (.A(_0867_),
    .B(_3115_),
    .Y(_1752_));
 sky130_fd_sc_hd__nand2_1 _5043_ (.A(_1751_),
    .B(_1752_),
    .Y(_1753_));
 sky130_fd_sc_hd__a221oi_2 _5044_ (.A1(_0385_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .C1(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__nand2_1 _5045_ (.A(_0874_),
    .B(_2904_),
    .Y(_1755_));
 sky130_fd_sc_hd__nand2_1 _5046_ (.A(_0877_),
    .B(_0346_),
    .Y(_1756_));
 sky130_fd_sc_hd__nand2_1 _5047_ (.A(_1755_),
    .B(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__a221oi_1 _5048_ (.A1(_0443_),
    .A2(_0872_),
    .B1(_0587_),
    .B2(_0873_),
    .C1(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__nand2_1 _5049_ (.A(_0895_),
    .B(_1011_),
    .Y(_1759_));
 sky130_fd_sc_hd__nand2_1 _5050_ (.A(_0897_),
    .B(_0894_),
    .Y(_1760_));
 sky130_fd_sc_hd__nand2_1 _5051_ (.A(_1759_),
    .B(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__a221oi_1 _5052_ (.A1(_0892_),
    .A2(_0464_),
    .B1(_0893_),
    .B2(_0742_),
    .C1(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__nand2_1 _5053_ (.A(_0883_),
    .B(_2881_),
    .Y(_1763_));
 sky130_fd_sc_hd__nand2_1 _5054_ (.A(_0885_),
    .B(_0551_),
    .Y(_1764_));
 sky130_fd_sc_hd__or2b_1 _5055_ (.A(_0889_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[71] ),
    .X(_1765_));
 sky130_fd_sc_hd__o2111a_1 _5056_ (.A1(_0984_),
    .A2(_0882_),
    .B1(_1763_),
    .C1(_1764_),
    .D1(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__and4_1 _5057_ (.A(_1754_),
    .B(_1758_),
    .C(_1762_),
    .D(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__and4_1 _5058_ (.A(_1724_),
    .B(_1738_),
    .C(_1750_),
    .D(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__o22ai_1 _5059_ (.A1(_1185_),
    .A2(_3131_),
    .B1(_3108_),
    .B2(_3135_),
    .Y(_1769_));
 sky130_fd_sc_hd__a221oi_1 _5060_ (.A1(_0336_),
    .A2(_3126_),
    .B1(_3146_),
    .B2(_3123_),
    .C1(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__nand2_1 _5061_ (.A(_3118_),
    .B(_0392_),
    .Y(_1771_));
 sky130_fd_sc_hd__o21ai_1 _5062_ (.A1(_1066_),
    .A2(_3110_),
    .B1(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__a221oi_1 _5063_ (.A1(_2951_),
    .A2(_0907_),
    .B1(_2957_),
    .B2(_0908_),
    .C1(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__nand2_1 _5064_ (.A(_3100_),
    .B(_0406_),
    .Y(_1774_));
 sky130_fd_sc_hd__o21ai_1 _5065_ (.A1(_0334_),
    .A2(_3093_),
    .B1(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__a221oi_2 _5066_ (.A1(_2974_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_0657_),
    .C1(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__or2_1 _5067_ (.A(_0602_),
    .B(_3080_),
    .X(_1777_));
 sky130_fd_sc_hd__or2_1 _5068_ (.A(_3011_),
    .B(_3084_),
    .X(_1778_));
 sky130_fd_sc_hd__nand2_1 _5069_ (.A(_3087_),
    .B(_3139_),
    .Y(_1779_));
 sky130_fd_sc_hd__o2111a_1 _5070_ (.A1(_0653_),
    .A2(_3077_),
    .B1(_1777_),
    .C1(_1778_),
    .D1(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__and4_1 _5071_ (.A(_1770_),
    .B(_1773_),
    .C(_1776_),
    .D(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__o22ai_1 _5072_ (.A1(_1017_),
    .A2(_0956_),
    .B1(_1256_),
    .B2(_0958_),
    .Y(_1782_));
 sky130_fd_sc_hd__a221oi_2 _5073_ (.A1(_2818_),
    .A2(_0954_),
    .B1(_2816_),
    .B2(_0955_),
    .C1(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__o22ai_1 _5074_ (.A1(_0730_),
    .A2(_0963_),
    .B1(_0543_),
    .B2(_0964_),
    .Y(_1784_));
 sky130_fd_sc_hd__a221oi_1 _5075_ (.A1(_2859_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_0709_),
    .C1(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__o22ai_1 _5076_ (.A1(_1075_),
    .A2(_0969_),
    .B1(_3129_),
    .B2(_0971_),
    .Y(_1786_));
 sky130_fd_sc_hd__a221oi_1 _5077_ (.A1(_0967_),
    .A2(_1116_),
    .B1(_0968_),
    .B2(_0841_),
    .C1(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__o22ai_1 _5078_ (.A1(_0574_),
    .A2(_0976_),
    .B1(_3075_),
    .B2(_0977_),
    .Y(_1788_));
 sky130_fd_sc_hd__a221oi_1 _5079_ (.A1(_0974_),
    .A2(_2939_),
    .B1(_0975_),
    .B2(_2926_),
    .C1(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__and4_1 _5080_ (.A(_1783_),
    .B(_1785_),
    .C(_1787_),
    .D(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__o22ai_1 _5081_ (.A1(_0641_),
    .A2(_0405_),
    .B1(_0506_),
    .B2(_0409_),
    .Y(_1791_));
 sky130_fd_sc_hd__a221oi_1 _5082_ (.A1(_0981_),
    .A2(_0402_),
    .B1(_0982_),
    .B2(_2863_),
    .C1(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_0990_),
    .B(_3002_),
    .Y(_1793_));
 sky130_fd_sc_hd__nand2_1 _5084_ (.A(_0992_),
    .B(_2990_),
    .Y(_1794_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_1793_),
    .B(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__a221oi_1 _5086_ (.A1(_2993_),
    .A2(_0987_),
    .B1(_0412_),
    .B2(_0989_),
    .C1(_1795_),
    .Y(_1796_));
 sky130_fd_sc_hd__nand2_1 _5087_ (.A(_0428_),
    .B(_0920_),
    .Y(_1797_));
 sky130_fd_sc_hd__nand2_1 _5088_ (.A(_0999_),
    .B(_0583_),
    .Y(_1798_));
 sky130_fd_sc_hd__nand2_1 _5089_ (.A(_1797_),
    .B(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__a221oi_1 _5090_ (.A1(_2848_),
    .A2(_0996_),
    .B1(_0495_),
    .B2(_0997_),
    .C1(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__a22o_1 _5091_ (.A1(_0439_),
    .A2(_3034_),
    .B1(_0441_),
    .B2(_3048_),
    .X(_1801_));
 sky130_fd_sc_hd__o22ai_1 _5092_ (.A1(_3067_),
    .A2(_0446_),
    .B1(_3031_),
    .B2(_0449_),
    .Y(_1802_));
 sky130_fd_sc_hd__nor2_1 _5093_ (.A(_1801_),
    .B(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__and4_1 _5094_ (.A(_1792_),
    .B(_1796_),
    .C(_1800_),
    .D(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__nand2_1 _5095_ (.A(_0925_),
    .B(_0420_),
    .Y(_1805_));
 sky130_fd_sc_hd__o21ai_1 _5096_ (.A1(_2849_),
    .A2(_0923_),
    .B1(_1805_),
    .Y(_1806_));
 sky130_fd_sc_hd__a221oi_1 _5097_ (.A1(_2987_),
    .A2(_0922_),
    .B1(_0607_),
    .B2(_0921_),
    .C1(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__nand2_1 _5098_ (.A(_0947_),
    .B(_0435_),
    .Y(_1808_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_0949_),
    .B(_0371_),
    .Y(_1809_));
 sky130_fd_sc_hd__nand2_1 _5100_ (.A(_1808_),
    .B(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__a221oi_1 _5101_ (.A1(_1000_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_2931_),
    .C1(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(_0939_),
    .B(_3132_),
    .Y(_1812_));
 sky130_fd_sc_hd__nand2_1 _5103_ (.A(_0941_),
    .B(_2830_),
    .Y(_1813_));
 sky130_fd_sc_hd__nand2_1 _5104_ (.A(_1812_),
    .B(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__a221oi_1 _5105_ (.A1(_0937_),
    .A2(_0656_),
    .B1(_0553_),
    .B2(_0938_),
    .C1(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__a22o_1 _5106_ (.A1(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .X(_1816_));
 sky130_fd_sc_hd__a22o_1 _5107_ (.A1(_0933_),
    .A2(_0638_),
    .B1(_0934_),
    .B2(_0610_),
    .X(_1817_));
 sky130_fd_sc_hd__nor2_1 _5108_ (.A(_1816_),
    .B(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__and4_1 _5109_ (.A(_1807_),
    .B(_1811_),
    .C(_1815_),
    .D(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__and4_1 _5110_ (.A(_1781_),
    .B(_1790_),
    .C(_1804_),
    .D(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__nand3_1 _5111_ (.A(_1768_),
    .B(_0903_),
    .C(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__o21a_1 _5112_ (.A1(_3101_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1822_));
 sky130_fd_sc_hd__nand2_1 _5113_ (.A(_1821_),
    .B(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__nand2_1 _5114_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_1824_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_1823_),
    .B(_1824_),
    .Y(_0294_));
 sky130_fd_sc_hd__a22o_1 _5116_ (.A1(\egd_top.BitStream_buffer.BS_buffer[6] ),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0988_),
    .X(_1825_));
 sky130_fd_sc_hd__a221oi_2 _5117_ (.A1(_2791_),
    .A2(_0782_),
    .B1(_1116_),
    .B2(_0781_),
    .C1(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__nand2_1 _5118_ (.A(_0791_),
    .B(_0330_),
    .Y(_1827_));
 sky130_fd_sc_hd__o21ai_1 _5119_ (.A1(_0538_),
    .A2(_0790_),
    .B1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__a221oi_1 _5120_ (.A1(_2804_),
    .A2(_0787_),
    .B1(_2907_),
    .B2(_0788_),
    .C1(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__nand2_1 _5121_ (.A(_0797_),
    .B(_2816_),
    .Y(_1830_));
 sky130_fd_sc_hd__o21ai_1 _5122_ (.A1(_1256_),
    .A2(_0796_),
    .B1(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__a31oi_1 _5123_ (.A1(_2822_),
    .A2(_2996_),
    .A3(_2927_),
    .B1(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5124_ (.A(_0802_),
    .B(_2810_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _5125_ (.A(_0804_),
    .B(_1011_),
    .Y(_1834_));
 sky130_fd_sc_hd__nand2_1 _5126_ (.A(_1833_),
    .B(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__a221oi_1 _5127_ (.A1(_2806_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_2828_),
    .C1(_1835_),
    .Y(_1836_));
 sky130_fd_sc_hd__and4_2 _5128_ (.A(_1826_),
    .B(_1829_),
    .C(_1832_),
    .D(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__nand2_1 _5129_ (.A(_0812_),
    .B(_2980_),
    .Y(_1838_));
 sky130_fd_sc_hd__o21ai_1 _5130_ (.A1(_1519_),
    .A2(_0811_),
    .B1(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__a221oi_1 _5131_ (.A1(_2808_),
    .A2(_0810_),
    .B1(_3070_),
    .B2(_0809_),
    .C1(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__nand2_1 _5132_ (.A(_0818_),
    .B(_0625_),
    .Y(_1841_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(_0820_),
    .B(_2826_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _5134_ (.A(_1841_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__a221oi_1 _5135_ (.A1(_0816_),
    .A2(_2800_),
    .B1(_0817_),
    .B2(_0777_),
    .C1(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__o22ai_1 _5136_ (.A1(_2914_),
    .A2(_0826_),
    .B1(_0506_),
    .B2(_0827_),
    .Y(_1845_));
 sky130_fd_sc_hd__a221oi_1 _5137_ (.A1(_0824_),
    .A2(_3127_),
    .B1(_0825_),
    .B2(_3124_),
    .C1(_1845_),
    .Y(_1846_));
 sky130_fd_sc_hd__nand2_1 _5138_ (.A(_0833_),
    .B(_2824_),
    .Y(_1847_));
 sky130_fd_sc_hd__nand2_1 _5139_ (.A(_0835_),
    .B(_2874_),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _5140_ (.A(_1847_),
    .B(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__a221oi_1 _5141_ (.A1(_0420_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_0458_),
    .C1(_1849_),
    .Y(_1850_));
 sky130_fd_sc_hd__and4_1 _5142_ (.A(_1840_),
    .B(_1844_),
    .C(_1846_),
    .D(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__nand2_1 _5143_ (.A(_0844_),
    .B(_3053_),
    .Y(_1852_));
 sky130_fd_sc_hd__o21ai_1 _5144_ (.A1(_0516_),
    .A2(_0843_),
    .B1(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__a221oi_1 _5145_ (.A1(_0412_),
    .A2(_0840_),
    .B1(_3007_),
    .B2(_0842_),
    .C1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__nand2_1 _5146_ (.A(_2867_),
    .B(_2935_),
    .Y(_1855_));
 sky130_fd_sc_hd__o21ai_1 _5147_ (.A1(_0881_),
    .A2(_0850_),
    .B1(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__a221oi_1 _5148_ (.A1(_3017_),
    .A2(_0848_),
    .B1(_2922_),
    .B2(_0849_),
    .C1(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_2858_),
    .B(_0926_),
    .Y(_1858_));
 sky130_fd_sc_hd__o21ai_1 _5150_ (.A1(_0789_),
    .A2(_2854_),
    .B1(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__a221oi_1 _5151_ (.A1(_0920_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0587_),
    .C1(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__o22ai_1 _5152_ (.A1(_0337_),
    .A2(_2912_),
    .B1(_1403_),
    .B2(_2917_),
    .Y(_1861_));
 sky130_fd_sc_hd__a221oi_1 _5153_ (.A1(_0378_),
    .A2(_0857_),
    .B1(_0341_),
    .B2(_0858_),
    .C1(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__and4_1 _5154_ (.A(_1854_),
    .B(_1857_),
    .C(_1860_),
    .D(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_0865_),
    .B(_2931_),
    .Y(_1864_));
 sky130_fd_sc_hd__nand2_1 _5156_ (.A(_0867_),
    .B(_0385_),
    .Y(_1865_));
 sky130_fd_sc_hd__nand2_1 _5157_ (.A(_1864_),
    .B(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__a221oi_1 _5158_ (.A1(_0389_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_3115_),
    .C1(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_0874_),
    .B(_0477_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand2_1 _5160_ (.A(_0877_),
    .B(_3112_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _5161_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__a221oi_1 _5162_ (.A1(_2987_),
    .A2(_0872_),
    .B1(_0742_),
    .B2(_0873_),
    .C1(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__nand2_1 _5163_ (.A(_0895_),
    .B(_0886_),
    .Y(_1872_));
 sky130_fd_sc_hd__nand2_1 _5164_ (.A(_0897_),
    .B(_1000_),
    .Y(_1873_));
 sky130_fd_sc_hd__nand2_1 _5165_ (.A(_1872_),
    .B(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__a221oi_1 _5166_ (.A1(_0892_),
    .A2(_2959_),
    .B1(_0893_),
    .B2(_0583_),
    .C1(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__nand2_1 _5167_ (.A(_0883_),
    .B(_2943_),
    .Y(_1876_));
 sky130_fd_sc_hd__nand2_1 _5168_ (.A(_0885_),
    .B(_2881_),
    .Y(_1877_));
 sky130_fd_sc_hd__or2b_1 _5169_ (.A(_0889_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[72] ),
    .X(_1878_));
 sky130_fd_sc_hd__o2111a_1 _5170_ (.A1(_0403_),
    .A2(_0882_),
    .B1(_1876_),
    .C1(_1877_),
    .D1(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__and4_1 _5171_ (.A(_1867_),
    .B(_1871_),
    .C(_1875_),
    .D(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__and4_1 _5172_ (.A(_1837_),
    .B(_1851_),
    .C(_1863_),
    .D(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__o22ai_1 _5173_ (.A1(_1301_),
    .A2(_3131_),
    .B1(_3129_),
    .B2(_3135_),
    .Y(_1882_));
 sky130_fd_sc_hd__a221oi_1 _5174_ (.A1(_3146_),
    .A2(_3126_),
    .B1(_3132_),
    .B2(_3123_),
    .C1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__nand2_1 _5175_ (.A(_3118_),
    .B(_3142_),
    .Y(_1884_));
 sky130_fd_sc_hd__o21ai_1 _5176_ (.A1(_1185_),
    .A2(_3110_),
    .B1(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__a221oi_1 _5177_ (.A1(_0392_),
    .A2(_0907_),
    .B1(_0371_),
    .B2(_0908_),
    .C1(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(_3100_),
    .B(_3040_),
    .Y(_1887_));
 sky130_fd_sc_hd__o21ai_1 _5179_ (.A1(_3144_),
    .A2(_3093_),
    .B1(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__a221oi_1 _5180_ (.A1(_0333_),
    .A2(_3096_),
    .B1(_3104_),
    .B2(_0894_),
    .C1(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__or2_1 _5181_ (.A(_0757_),
    .B(_3080_),
    .X(_1890_));
 sky130_fd_sc_hd__or2_1 _5182_ (.A(_0407_),
    .B(_3084_),
    .X(_1891_));
 sky130_fd_sc_hd__nand2_1 _5183_ (.A(_3087_),
    .B(_0398_),
    .Y(_1892_));
 sky130_fd_sc_hd__o2111a_1 _5184_ (.A1(_0888_),
    .A2(_3077_),
    .B1(_1890_),
    .C1(_1891_),
    .D1(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__and4_1 _5185_ (.A(_1883_),
    .B(_1886_),
    .C(_1889_),
    .D(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__o22ai_2 _5186_ (.A1(_3067_),
    .A2(_0956_),
    .B1(_1372_),
    .B2(_0958_),
    .Y(_1895_));
 sky130_fd_sc_hd__a221oi_4 _5187_ (.A1(_2820_),
    .A2(_0954_),
    .B1(_2818_),
    .B2(_0955_),
    .C1(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__o22ai_1 _5188_ (.A1(_3075_),
    .A2(_0963_),
    .B1(_3108_),
    .B2(_0964_),
    .Y(_1897_));
 sky130_fd_sc_hd__a221oi_1 _5189_ (.A1(_2830_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_2859_),
    .C1(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__o22ai_1 _5190_ (.A1(_2952_),
    .A2(_0969_),
    .B1(_0561_),
    .B2(_0971_),
    .Y(_1899_));
 sky130_fd_sc_hd__a221oi_1 _5191_ (.A1(_0967_),
    .A2(_0841_),
    .B1(_0968_),
    .B2(_3101_),
    .C1(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__o22ai_1 _5192_ (.A1(_0730_),
    .A2(_0976_),
    .B1(_0543_),
    .B2(_0977_),
    .Y(_1901_));
 sky130_fd_sc_hd__a221oi_1 _5193_ (.A1(_0974_),
    .A2(_2926_),
    .B1(_0975_),
    .B2(_0346_),
    .C1(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hd__and4_1 _5194_ (.A(_1896_),
    .B(_1898_),
    .C(_1900_),
    .D(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__o22ai_1 _5195_ (.A1(_0859_),
    .A2(_0405_),
    .B1(_3091_),
    .B2(_0409_),
    .Y(_1904_));
 sky130_fd_sc_hd__a221oi_1 _5196_ (.A1(_0981_),
    .A2(_2863_),
    .B1(_0982_),
    .B2(_2920_),
    .C1(_1904_),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _5197_ (.A(_0990_),
    .B(_3030_),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _5198_ (.A(_0992_),
    .B(_3058_),
    .Y(_1907_));
 sky130_fd_sc_hd__nand2_1 _5199_ (.A(_1906_),
    .B(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__a221oi_1 _5200_ (.A1(_3010_),
    .A2(_0987_),
    .B1(_0414_),
    .B2(_0989_),
    .C1(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__nand2_1 _5201_ (.A(_0428_),
    .B(_0875_),
    .Y(_1910_));
 sky130_fd_sc_hd__nand2_1 _5202_ (.A(_0999_),
    .B(_0871_),
    .Y(_1911_));
 sky130_fd_sc_hd__nand2_1 _5203_ (.A(_1910_),
    .B(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__a221oi_1 _5204_ (.A1(_0464_),
    .A2(_0996_),
    .B1(_0657_),
    .B2(_0997_),
    .C1(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__a22o_1 _5205_ (.A1(_0439_),
    .A2(_3048_),
    .B1(_0441_),
    .B2(_3002_),
    .X(_1914_));
 sky130_fd_sc_hd__o22ai_1 _5206_ (.A1(_3154_),
    .A2(_0446_),
    .B1(_0526_),
    .B2(_0449_),
    .Y(_1915_));
 sky130_fd_sc_hd__nor2_1 _5207_ (.A(_1914_),
    .B(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hd__and4_1 _5208_ (.A(_1905_),
    .B(_1909_),
    .C(_1913_),
    .D(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__nand2_1 _5209_ (.A(_0925_),
    .B(_0607_),
    .Y(_1918_));
 sky130_fd_sc_hd__o21ai_1 _5210_ (.A1(_0465_),
    .A2(_0923_),
    .B1(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__a221oi_1 _5211_ (.A1(_3034_),
    .A2(_0922_),
    .B1(_2904_),
    .B2(_0921_),
    .C1(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__nand2_1 _5212_ (.A(_0947_),
    .B(_2957_),
    .Y(_1921_));
 sky130_fd_sc_hd__nand2_1 _5213_ (.A(_0949_),
    .B(_0656_),
    .Y(_1922_));
 sky130_fd_sc_hd__nand2_1 _5214_ (.A(_1921_),
    .B(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__a221oi_1 _5215_ (.A1(_0830_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_2939_),
    .C1(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_0939_),
    .B(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .Y(_1925_));
 sky130_fd_sc_hd__nand2_1 _5217_ (.A(_0941_),
    .B(\egd_top.BitStream_buffer.BS_buffer[76] ),
    .Y(_1926_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(_1925_),
    .B(_1926_),
    .Y(_1927_));
 sky130_fd_sc_hd__a221oi_1 _5219_ (.A1(_0937_),
    .A2(_3105_),
    .B1(_0709_),
    .B2(_0938_),
    .C1(_1927_),
    .Y(_1928_));
 sky130_fd_sc_hd__a22o_1 _5220_ (.A1(\egd_top.BitStream_buffer.BS_buffer[77] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .X(_1929_));
 sky130_fd_sc_hd__a22o_1 _5221_ (.A1(_0933_),
    .A2(_0610_),
    .B1(_0934_),
    .B2(_0443_),
    .X(_1930_));
 sky130_fd_sc_hd__nor2_1 _5222_ (.A(_1929_),
    .B(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__and4_1 _5223_ (.A(_1920_),
    .B(_1924_),
    .C(_1928_),
    .D(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__and4_1 _5224_ (.A(_1894_),
    .B(_1903_),
    .C(_1917_),
    .D(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__nand3_1 _5225_ (.A(_1881_),
    .B(_0903_),
    .C(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hd__o21a_1 _5226_ (.A1(_0551_),
    .A2(_0457_),
    .B1(_2790_),
    .X(_1935_));
 sky130_fd_sc_hd__nand2_1 _5227_ (.A(_1934_),
    .B(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _5228_ (.A(_0461_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _5229_ (.A(_1936_),
    .B(_1937_),
    .Y(_0293_));
 sky130_fd_sc_hd__a22o_1 _5230_ (.A1(_0988_),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_1116_),
    .X(_1938_));
 sky130_fd_sc_hd__a221oi_1 _5231_ (.A1(_2800_),
    .A2(_0782_),
    .B1(_0841_),
    .B2(_0781_),
    .C1(_1938_),
    .Y(_1939_));
 sky130_fd_sc_hd__nand2_1 _5232_ (.A(_0791_),
    .B(_2791_),
    .Y(_1940_));
 sky130_fd_sc_hd__o21ai_1 _5233_ (.A1(_0698_),
    .A2(_0790_),
    .B1(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__a221oi_1 _5234_ (.A1(_2806_),
    .A2(_0787_),
    .B1(_3127_),
    .B2(_0788_),
    .C1(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5235_ (.A(_0797_),
    .B(_2818_),
    .Y(_1943_));
 sky130_fd_sc_hd__o21ai_1 _5236_ (.A1(_1372_),
    .A2(_0796_),
    .B1(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__a31oi_1 _5237_ (.A1(_2824_),
    .A2(_2996_),
    .A3(_2927_),
    .B1(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__nand2_1 _5238_ (.A(_0802_),
    .B(_2812_),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(_0804_),
    .B(_0886_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _5240_ (.A(_1946_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__a221oi_1 _5241_ (.A1(_2808_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_0458_),
    .C1(_1948_),
    .Y(_1949_));
 sky130_fd_sc_hd__and4_2 _5242_ (.A(_1939_),
    .B(_1942_),
    .C(_1945_),
    .D(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_0812_),
    .B(_3097_),
    .Y(_1951_));
 sky130_fd_sc_hd__o21ai_1 _5244_ (.A1(_0334_),
    .A2(_0811_),
    .B1(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__a221oi_1 _5245_ (.A1(_2810_),
    .A2(_0810_),
    .B1(_0330_),
    .B2(_0809_),
    .C1(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__nand2_1 _5246_ (.A(_0818_),
    .B(_0777_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(_0820_),
    .B(_2828_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand2_1 _5248_ (.A(_1954_),
    .B(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__a221oi_2 _5249_ (.A1(_0816_),
    .A2(_2802_),
    .B1(_0817_),
    .B2(_1011_),
    .C1(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__o22ai_1 _5250_ (.A1(_2981_),
    .A2(_0826_),
    .B1(_3091_),
    .B2(_0827_),
    .Y(_1958_));
 sky130_fd_sc_hd__a221oi_1 _5251_ (.A1(_0824_),
    .A2(_3124_),
    .B1(_0825_),
    .B2(_0395_),
    .C1(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(_0833_),
    .B(_2826_),
    .Y(_1960_));
 sky130_fd_sc_hd__nand2_1 _5253_ (.A(_0835_),
    .B(_0469_),
    .Y(_1961_));
 sky130_fd_sc_hd__nand2_1 _5254_ (.A(_1960_),
    .B(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__a221oi_1 _5255_ (.A1(_0607_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_0625_),
    .C1(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__and4_1 _5256_ (.A(_1953_),
    .B(_1957_),
    .C(_1959_),
    .D(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__nand2_1 _5257_ (.A(_0844_),
    .B(_2990_),
    .Y(_1965_));
 sky130_fd_sc_hd__o21ai_1 _5258_ (.A1(_3011_),
    .A2(_0843_),
    .B1(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__a221oi_1 _5259_ (.A1(_0414_),
    .A2(_0840_),
    .B1(_2993_),
    .B2(_0842_),
    .C1(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__nand2_1 _5260_ (.A(_2867_),
    .B(_0378_),
    .Y(_1968_));
 sky130_fd_sc_hd__o21ai_1 _5261_ (.A1(_3008_),
    .A2(_0850_),
    .B1(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__a221oi_1 _5262_ (.A1(_0402_),
    .A2(_0848_),
    .B1(_2913_),
    .B2(_0849_),
    .C1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand2_1 _5263_ (.A(_2858_),
    .B(_0920_),
    .Y(_1971_));
 sky130_fd_sc_hd__o21ai_1 _5264_ (.A1(_1017_),
    .A2(_2854_),
    .B1(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__a221oi_1 _5265_ (.A1(_0875_),
    .A2(_2840_),
    .B1(_2847_),
    .B2(_0742_),
    .C1(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__o22ai_1 _5266_ (.A1(_3147_),
    .A2(_2911_),
    .B1(_1519_),
    .B2(_2916_),
    .Y(_1974_));
 sky130_fd_sc_hd__a221oi_1 _5267_ (.A1(_0341_),
    .A2(_0857_),
    .B1(_0343_),
    .B2(_0858_),
    .C1(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__and4_1 _5268_ (.A(_1967_),
    .B(_1970_),
    .C(_1973_),
    .D(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__nand2_1 _5269_ (.A(_0865_),
    .B(_2939_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _5270_ (.A(_0867_),
    .B(_0389_),
    .Y(_1978_));
 sky130_fd_sc_hd__nand2_1 _5271_ (.A(_1977_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__a221oi_2 _5272_ (.A1(_2951_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_0385_),
    .C1(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__nand2_1 _5273_ (.A(_0874_),
    .B(_0638_),
    .Y(_1981_));
 sky130_fd_sc_hd__nand2_1 _5274_ (.A(_0877_),
    .B(_3119_),
    .Y(_1982_));
 sky130_fd_sc_hd__nand2_1 _5275_ (.A(_1981_),
    .B(_1982_),
    .Y(_1983_));
 sky130_fd_sc_hd__a221oi_1 _5276_ (.A1(_3034_),
    .A2(_0872_),
    .B1(_0583_),
    .B2(_0873_),
    .C1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__nand2_1 _5277_ (.A(_0895_),
    .B(_2874_),
    .Y(_1985_));
 sky130_fd_sc_hd__nand2_1 _5278_ (.A(_0897_),
    .B(_0830_),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_1 _5279_ (.A(_1985_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__a221oi_1 _5280_ (.A1(_0892_),
    .A2(_0495_),
    .B1(_0893_),
    .B2(_0871_),
    .C1(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5281_ (.A(_0883_),
    .B(_0412_),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _5282_ (.A(_0885_),
    .B(_2943_),
    .Y(_1990_));
 sky130_fd_sc_hd__or2b_1 _5283_ (.A(_0889_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[73] ),
    .X(_1991_));
 sky130_fd_sc_hd__o2111a_1 _5284_ (.A1(_0601_),
    .A2(_0882_),
    .B1(_1989_),
    .C1(_1990_),
    .D1(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__and4_1 _5285_ (.A(_1980_),
    .B(_1984_),
    .C(_1988_),
    .D(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__and4_1 _5286_ (.A(_1950_),
    .B(_1964_),
    .C(_1976_),
    .D(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__o22ai_1 _5287_ (.A1(_1052_),
    .A2(_0404_),
    .B1(_2908_),
    .B2(_0408_),
    .Y(_1995_));
 sky130_fd_sc_hd__a221oi_1 _5288_ (.A1(_0981_),
    .A2(_2920_),
    .B1(_0982_),
    .B2(_2922_),
    .C1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_1 _5289_ (.A(_0990_),
    .B(_3037_),
    .Y(_1997_));
 sky130_fd_sc_hd__nand2_1 _5290_ (.A(_0992_),
    .B(_3066_),
    .Y(_1998_));
 sky130_fd_sc_hd__nand2_1 _5291_ (.A(_1997_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__a221oi_1 _5292_ (.A1(_0406_),
    .A2(_0987_),
    .B1(_2887_),
    .B2(_0989_),
    .C1(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__nand2_1 _5293_ (.A(_0427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[88] ),
    .Y(_2001_));
 sky130_fd_sc_hd__nand2_1 _5294_ (.A(_0999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[92] ),
    .Y(_2002_));
 sky130_fd_sc_hd__nand2_1 _5295_ (.A(_2001_),
    .B(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__a221oi_2 _5296_ (.A1(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .A2(_0996_),
    .B1(\egd_top.BitStream_buffer.BS_buffer[82] ),
    .B2(_0997_),
    .C1(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__a22o_1 _5297_ (.A1(_0438_),
    .A2(_3002_),
    .B1(_0440_),
    .B2(_3030_),
    .X(_2005_));
 sky130_fd_sc_hd__o22ai_1 _5298_ (.A1(_0567_),
    .A2(_0445_),
    .B1(_0686_),
    .B2(_0448_),
    .Y(_2006_));
 sky130_fd_sc_hd__nor2_1 _5299_ (.A(_2005_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__and4_1 _5300_ (.A(_1996_),
    .B(_2000_),
    .C(_2004_),
    .D(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__nand2_1 _5301_ (.A(_3117_),
    .B(_3139_),
    .Y(_2009_));
 sky130_fd_sc_hd__o21ai_1 _5302_ (.A1(_1301_),
    .A2(_3109_),
    .B1(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__a221oi_1 _5303_ (.A1(_3142_),
    .A2(_0907_),
    .B1(_0656_),
    .B2(_0908_),
    .C1(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _5304_ (.A(_3099_),
    .B(_3015_),
    .Y(_2012_));
 sky130_fd_sc_hd__o21ai_1 _5305_ (.A1(_0337_),
    .A2(_3092_),
    .B1(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hd__a221oi_2 _5306_ (.A1(_3143_),
    .A2(_3095_),
    .B1(_3103_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[83] ),
    .C1(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__or2_1 _5307_ (.A(_0984_),
    .B(_3079_),
    .X(_2015_));
 sky130_fd_sc_hd__or2_1 _5308_ (.A(_0602_),
    .B(_3083_),
    .X(_2016_));
 sky130_fd_sc_hd__nand2_1 _5309_ (.A(_3086_),
    .B(_0366_),
    .Y(_2017_));
 sky130_fd_sc_hd__o2111a_1 _5310_ (.A1(_1066_),
    .A2(_3076_),
    .B1(_2015_),
    .C1(_2016_),
    .D1(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__a22o_1 _5311_ (.A1(_3122_),
    .A2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .B1(_3125_),
    .B2(_3132_),
    .X(_2019_));
 sky130_fd_sc_hd__o22ai_1 _5312_ (.A1(_1417_),
    .A2(_3130_),
    .B1(_0561_),
    .B2(_3134_),
    .Y(_2020_));
 sky130_fd_sc_hd__nor2_1 _5313_ (.A(_2019_),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__and4_1 _5314_ (.A(_2011_),
    .B(_2014_),
    .C(_2018_),
    .D(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__and2_1 _5315_ (.A(_2008_),
    .B(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__a22o_1 _5316_ (.A1(\egd_top.BitStream_buffer.BS_buffer[78] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_0657_),
    .X(_2024_));
 sky130_fd_sc_hd__a221oi_1 _5317_ (.A1(_0443_),
    .A2(_0933_),
    .B1(_2987_),
    .B2(_0934_),
    .C1(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _5318_ (.A(_0925_),
    .B(_2904_),
    .Y(_2026_));
 sky130_fd_sc_hd__o21ai_1 _5319_ (.A1(_3151_),
    .A2(_0923_),
    .B1(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__a221oi_1 _5320_ (.A1(_3048_),
    .A2(_0922_),
    .B1(_0477_),
    .B2(_0921_),
    .C1(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _5321_ (.A(_0939_),
    .B(_2931_),
    .Y(_2029_));
 sky130_fd_sc_hd__nand2_1 _5322_ (.A(_0941_),
    .B(_2848_),
    .Y(_2030_));
 sky130_fd_sc_hd__nand2_1 _5323_ (.A(_2029_),
    .B(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__a221oi_1 _5324_ (.A1(_0937_),
    .A2(_0553_),
    .B1(_2859_),
    .B2(_0938_),
    .C1(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(_0947_),
    .B(_0371_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand2_1 _5326_ (.A(_0949_),
    .B(_3105_),
    .Y(_2034_));
 sky130_fd_sc_hd__nand2_1 _5327_ (.A(_2033_),
    .B(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__a221oi_1 _5328_ (.A1(_0926_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_2926_),
    .C1(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__and4_1 _5329_ (.A(_2025_),
    .B(_2028_),
    .C(_2032_),
    .D(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__o22ai_2 _5330_ (.A1(_3154_),
    .A2(_0956_),
    .B1(_1488_),
    .B2(_0958_),
    .Y(_2038_));
 sky130_fd_sc_hd__a221oi_4 _5331_ (.A1(_2822_),
    .A2(_0954_),
    .B1(_2820_),
    .B2(_0955_),
    .C1(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__o22ai_1 _5332_ (.A1(_0543_),
    .A2(_0963_),
    .B1(_3129_),
    .B2(_0964_),
    .Y(_2040_));
 sky130_fd_sc_hd__a221oi_1 _5333_ (.A1(_0463_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_2830_),
    .C1(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__o22ai_1 _5334_ (.A1(_0492_),
    .A2(_0969_),
    .B1(_0717_),
    .B2(_0971_),
    .Y(_2042_));
 sky130_fd_sc_hd__a221oi_1 _5335_ (.A1(_0967_),
    .A2(_3101_),
    .B1(_0968_),
    .B2(_0551_),
    .C1(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__o22ai_1 _5336_ (.A1(_3075_),
    .A2(_0976_),
    .B1(_3108_),
    .B2(_0977_),
    .Y(_2044_));
 sky130_fd_sc_hd__a221oi_1 _5337_ (.A1(_0974_),
    .A2(_0346_),
    .B1(_0975_),
    .B2(_3112_),
    .C1(_2044_),
    .Y(_2045_));
 sky130_fd_sc_hd__and4_2 _5338_ (.A(_2039_),
    .B(_2041_),
    .C(_2043_),
    .D(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__and3_1 _5339_ (.A(_2023_),
    .B(_2037_),
    .C(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__nand3_1 _5340_ (.A(_1994_),
    .B(_0903_),
    .C(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__o21a_1 _5341_ (.A1(_2881_),
    .A2(_0456_),
    .B1(_2790_),
    .X(_2049_));
 sky130_fd_sc_hd__nand2_1 _5342_ (.A(_2048_),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__nand2_1 _5343_ (.A(net221),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2051_));
 sky130_fd_sc_hd__nand2_1 _5344_ (.A(_2050_),
    .B(_2051_),
    .Y(_0292_));
 sky130_fd_sc_hd__a22o_1 _5345_ (.A1(_1116_),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0841_),
    .X(_2052_));
 sky130_fd_sc_hd__a221oi_1 _5346_ (.A1(_2802_),
    .A2(_0782_),
    .B1(_3101_),
    .B2(_0781_),
    .C1(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _5347_ (.A(_0791_),
    .B(_2800_),
    .Y(_2054_));
 sky130_fd_sc_hd__o21ai_1 _5348_ (.A1(_0795_),
    .A2(_0790_),
    .B1(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__a221oi_1 _5349_ (.A1(_2808_),
    .A2(_0787_),
    .B1(_3124_),
    .B2(_0788_),
    .C1(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _5350_ (.A(_0797_),
    .B(_2820_),
    .Y(_2057_));
 sky130_fd_sc_hd__o21ai_1 _5351_ (.A1(_1488_),
    .A2(_0796_),
    .B1(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__a31oi_1 _5352_ (.A1(_2826_),
    .A2(_2996_),
    .A3(_2927_),
    .B1(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__nand2_1 _5353_ (.A(_0802_),
    .B(_2814_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _5354_ (.A(_0804_),
    .B(_2874_),
    .Y(_2061_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_2060_),
    .B(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__a221oi_1 _5356_ (.A1(_2810_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_0625_),
    .C1(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__and4_2 _5357_ (.A(_2053_),
    .B(_2056_),
    .C(_2059_),
    .D(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__nand2_1 _5358_ (.A(_0812_),
    .B(_3090_),
    .Y(_2065_));
 sky130_fd_sc_hd__o21ai_1 _5359_ (.A1(_3144_),
    .A2(_0811_),
    .B1(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__a221oi_1 _5360_ (.A1(_2791_),
    .A2(_0809_),
    .B1(_2812_),
    .B2(_0810_),
    .C1(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__nand2_1 _5361_ (.A(_0818_),
    .B(_1011_),
    .Y(_2068_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(_0820_),
    .B(_0458_),
    .Y(_2069_));
 sky130_fd_sc_hd__nand2_1 _5363_ (.A(_2068_),
    .B(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__a221oi_1 _5364_ (.A1(_0816_),
    .A2(_2804_),
    .B1(_0817_),
    .B2(_0886_),
    .C1(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hd__o22ai_1 _5365_ (.A1(_0506_),
    .A2(_0826_),
    .B1(_2908_),
    .B2(_0827_),
    .Y(_2072_));
 sky130_fd_sc_hd__a221oi_1 _5366_ (.A1(_0824_),
    .A2(_0395_),
    .B1(_0825_),
    .B2(_2935_),
    .C1(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__nand2_1 _5367_ (.A(_0833_),
    .B(_2828_),
    .Y(_2074_));
 sky130_fd_sc_hd__nand2_1 _5368_ (.A(_0835_),
    .B(_0988_),
    .Y(_2075_));
 sky130_fd_sc_hd__nand2_1 _5369_ (.A(_2074_),
    .B(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__a221oi_1 _5370_ (.A1(_2904_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_0777_),
    .C1(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__and4_1 _5371_ (.A(_2067_),
    .B(_2071_),
    .C(_2073_),
    .D(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__nand2_1 _5372_ (.A(_0844_),
    .B(_3058_),
    .Y(_2079_));
 sky130_fd_sc_hd__o21ai_1 _5373_ (.A1(_0407_),
    .A2(_0843_),
    .B1(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__a221oi_1 _5374_ (.A1(_2887_),
    .A2(_0840_),
    .B1(_3010_),
    .B2(_0842_),
    .C1(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_1 _5375_ (.A(_2866_),
    .B(_0341_),
    .Y(_2082_));
 sky130_fd_sc_hd__o21ai_1 _5376_ (.A1(_0516_),
    .A2(_0850_),
    .B1(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__a221oi_1 _5377_ (.A1(_2863_),
    .A2(_0848_),
    .B1(_2980_),
    .B2(_0849_),
    .C1(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(_2857_),
    .B(_0875_),
    .Y(_2085_));
 sky130_fd_sc_hd__o21ai_1 _5379_ (.A1(_3067_),
    .A2(_2853_),
    .B1(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__a221oi_1 _5380_ (.A1(_0587_),
    .A2(_2839_),
    .B1(_2846_),
    .B2(_0583_),
    .C1(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__o22ai_1 _5381_ (.A1(_3133_),
    .A2(_2911_),
    .B1(_0334_),
    .B2(_2916_),
    .Y(_2088_));
 sky130_fd_sc_hd__a221oi_2 _5382_ (.A1(_0343_),
    .A2(_0857_),
    .B1(_2974_),
    .B2(_0858_),
    .C1(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__and4_1 _5383_ (.A(_2081_),
    .B(_2084_),
    .C(_2087_),
    .D(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__nand2_1 _5384_ (.A(_0865_),
    .B(_2926_),
    .Y(_2091_));
 sky130_fd_sc_hd__nand2_1 _5385_ (.A(_0867_),
    .B(_2951_),
    .Y(_2092_));
 sky130_fd_sc_hd__nand2_1 _5386_ (.A(_2091_),
    .B(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__a221oi_2 _5387_ (.A1(_0392_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_0389_),
    .C1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__nand2_1 _5388_ (.A(_0874_),
    .B(_0610_),
    .Y(_2095_));
 sky130_fd_sc_hd__nand2_1 _5389_ (.A(_0877_),
    .B(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(_2095_),
    .B(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__a221oi_1 _5391_ (.A1(_3048_),
    .A2(_0872_),
    .B1(_0871_),
    .B2(_0873_),
    .C1(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__nand2_1 _5392_ (.A(_0895_),
    .B(_0469_),
    .Y(_2099_));
 sky130_fd_sc_hd__nand2_1 _5393_ (.A(_0897_),
    .B(_0926_),
    .Y(_2100_));
 sky130_fd_sc_hd__nand2_1 _5394_ (.A(_2099_),
    .B(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__a221oi_1 _5395_ (.A1(_0892_),
    .A2(_0657_),
    .B1(_0893_),
    .B2(_0420_),
    .C1(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand2_1 _5396_ (.A(_0883_),
    .B(_0414_),
    .Y(_2103_));
 sky130_fd_sc_hd__nand2_1 _5397_ (.A(_0885_),
    .B(_0412_),
    .Y(_2104_));
 sky130_fd_sc_hd__or2b_1 _5398_ (.A(_0889_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[74] ),
    .X(_2105_));
 sky130_fd_sc_hd__o2111a_1 _5399_ (.A1(_0756_),
    .A2(_0882_),
    .B1(_2103_),
    .C1(_2104_),
    .D1(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__and4_1 _5400_ (.A(_2094_),
    .B(_2098_),
    .C(_2102_),
    .D(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__and4_1 _5401_ (.A(_2064_),
    .B(_2078_),
    .C(_2090_),
    .D(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__o22ai_1 _5402_ (.A1(_1171_),
    .A2(_0404_),
    .B1(_0480_),
    .B2(_0408_),
    .Y(_2109_));
 sky130_fd_sc_hd__a221oi_1 _5403_ (.A1(_0981_),
    .A2(_2922_),
    .B1(_0982_),
    .B2(_2913_),
    .C1(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(_0990_),
    .B(_3053_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_1 _5405_ (.A(_0992_),
    .B(_3153_),
    .Y(_2112_));
 sky130_fd_sc_hd__nand2_1 _5406_ (.A(_2111_),
    .B(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__a221oi_1 _5407_ (.A1(_3040_),
    .A2(_0987_),
    .B1(_3007_),
    .B2(_0989_),
    .C1(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_0427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[89] ),
    .Y(_2115_));
 sky130_fd_sc_hd__nand2_1 _5409_ (.A(_0999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[93] ),
    .Y(_2116_));
 sky130_fd_sc_hd__nand2_1 _5410_ (.A(_2115_),
    .B(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__a221oi_1 _5411_ (.A1(\egd_top.BitStream_buffer.BS_buffer[80] ),
    .A2(_0996_),
    .B1(_1000_),
    .B2(_0997_),
    .C1(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__a22o_1 _5412_ (.A1(_0438_),
    .A2(_3030_),
    .B1(_0440_),
    .B2(_3037_),
    .X(_2119_));
 sky130_fd_sc_hd__o22ai_1 _5413_ (.A1(_0723_),
    .A2(_0445_),
    .B1(_0789_),
    .B2(_0448_),
    .Y(_2120_));
 sky130_fd_sc_hd__nor2_1 _5414_ (.A(_2119_),
    .B(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__and4_1 _5415_ (.A(_2110_),
    .B(_2114_),
    .C(_2118_),
    .D(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__nand2_1 _5416_ (.A(_3117_),
    .B(_0398_),
    .Y(_2123_));
 sky130_fd_sc_hd__o21ai_1 _5417_ (.A1(_1417_),
    .A2(_3109_),
    .B1(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__a221oi_1 _5418_ (.A1(_3139_),
    .A2(_0907_),
    .B1(_3105_),
    .B2(_0908_),
    .C1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__nand2_1 _5419_ (.A(_3099_),
    .B(_3017_),
    .Y(_2126_));
 sky130_fd_sc_hd__o21ai_1 _5420_ (.A1(_3147_),
    .A2(_3092_),
    .B1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__a221oi_2 _5421_ (.A1(_0336_),
    .A2(_3095_),
    .B1(_3103_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[84] ),
    .C1(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__or2_1 _5422_ (.A(_0403_),
    .B(_3079_),
    .X(_2129_));
 sky130_fd_sc_hd__or2_1 _5423_ (.A(_0757_),
    .B(_3083_),
    .X(_2130_));
 sky130_fd_sc_hd__nand2_1 _5424_ (.A(_3086_),
    .B(_0435_),
    .Y(_2131_));
 sky130_fd_sc_hd__o2111a_1 _5425_ (.A1(_1185_),
    .A2(_3076_),
    .B1(_2129_),
    .C1(_2130_),
    .D1(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__a22o_1 _5426_ (.A1(_3122_),
    .A2(_2931_),
    .B1(_3125_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .X(_2133_));
 sky130_fd_sc_hd__o22ai_1 _5427_ (.A1(_1533_),
    .A2(_3130_),
    .B1(_0717_),
    .B2(_3134_),
    .Y(_2134_));
 sky130_fd_sc_hd__nor2_1 _5428_ (.A(_2133_),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__and4_1 _5429_ (.A(_2125_),
    .B(_2128_),
    .C(_2132_),
    .D(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__and2_1 _5430_ (.A(_2122_),
    .B(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__a22o_1 _5431_ (.A1(\egd_top.BitStream_buffer.BS_buffer[79] ),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_0894_),
    .X(_2138_));
 sky130_fd_sc_hd__a221oi_1 _5432_ (.A1(_2987_),
    .A2(_0933_),
    .B1(_3034_),
    .B2(_0934_),
    .C1(_2138_),
    .Y(_2139_));
 sky130_fd_sc_hd__nand2_1 _5433_ (.A(_0925_),
    .B(_0477_),
    .Y(_2140_));
 sky130_fd_sc_hd__o21ai_1 _5434_ (.A1(_0444_),
    .A2(_0923_),
    .B1(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__a221oi_1 _5435_ (.A1(_0638_),
    .A2(_0921_),
    .B1(_3002_),
    .B2(_0922_),
    .C1(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(_0939_),
    .B(_2939_),
    .Y(_2143_));
 sky130_fd_sc_hd__nand2_1 _5437_ (.A(_0941_),
    .B(_0464_),
    .Y(_2144_));
 sky130_fd_sc_hd__nand2_1 _5438_ (.A(_2143_),
    .B(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__a221oi_1 _5439_ (.A1(_0937_),
    .A2(_0709_),
    .B1(_2830_),
    .B2(_0938_),
    .C1(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(_0947_),
    .B(_0656_),
    .Y(_2147_));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(_0949_),
    .B(_0553_),
    .Y(_2148_));
 sky130_fd_sc_hd__nand2_1 _5442_ (.A(_2147_),
    .B(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__a221oi_1 _5443_ (.A1(_0920_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_0346_),
    .C1(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__and4_1 _5444_ (.A(_2139_),
    .B(_2142_),
    .C(_2146_),
    .D(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__o22ai_1 _5445_ (.A1(_0567_),
    .A2(_0956_),
    .B1(_1603_),
    .B2(_0958_),
    .Y(_2152_));
 sky130_fd_sc_hd__a221oi_2 _5446_ (.A1(_2824_),
    .A2(_0954_),
    .B1(_2822_),
    .B2(_0955_),
    .C1(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__o22ai_1 _5447_ (.A1(_3108_),
    .A2(_0963_),
    .B1(_0561_),
    .B2(_0964_),
    .Y(_2154_));
 sky130_fd_sc_hd__a221oi_1 _5448_ (.A1(_2848_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_0463_),
    .C1(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__o22ai_1 _5449_ (.A1(_0653_),
    .A2(_0969_),
    .B1(_0904_),
    .B2(_0971_),
    .Y(_2156_));
 sky130_fd_sc_hd__a221oi_1 _5450_ (.A1(_0967_),
    .A2(_0551_),
    .B1(_0968_),
    .B2(_2881_),
    .C1(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__o22ai_1 _5451_ (.A1(_0543_),
    .A2(_0976_),
    .B1(_3129_),
    .B2(_0977_),
    .Y(_2158_));
 sky130_fd_sc_hd__a221oi_1 _5452_ (.A1(_0974_),
    .A2(_3112_),
    .B1(_0975_),
    .B2(_3119_),
    .C1(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__and4_1 _5453_ (.A(_2153_),
    .B(_2155_),
    .C(_2157_),
    .D(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__and3_1 _5454_ (.A(_2137_),
    .B(_2151_),
    .C(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__nand3_1 _5455_ (.A(_2108_),
    .B(_0903_),
    .C(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__o21a_1 _5456_ (.A1(_2943_),
    .A2(_0456_),
    .B1(_2790_),
    .X(_2163_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(_2162_),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(net221),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2165_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_2164_),
    .B(_2165_),
    .Y(_0291_));
 sky130_fd_sc_hd__a22o_1 _5460_ (.A1(_0841_),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_3101_),
    .X(_2166_));
 sky130_fd_sc_hd__a221oi_1 _5461_ (.A1(_2804_),
    .A2(_0782_),
    .B1(_0551_),
    .B2(_0781_),
    .C1(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__nand2_1 _5462_ (.A(_0791_),
    .B(_2802_),
    .Y(_2168_));
 sky130_fd_sc_hd__o21ai_1 _5463_ (.A1(_1021_),
    .A2(_0790_),
    .B1(_2168_),
    .Y(_2169_));
 sky130_fd_sc_hd__a221oi_1 _5464_ (.A1(_2810_),
    .A2(_0787_),
    .B1(_0395_),
    .B2(_0788_),
    .C1(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_0797_),
    .B(_2822_),
    .Y(_2171_));
 sky130_fd_sc_hd__o21ai_1 _5466_ (.A1(_1603_),
    .A2(_0796_),
    .B1(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__a31oi_1 _5467_ (.A1(_2828_),
    .A2(_2996_),
    .A3(_2927_),
    .B1(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__nand2_1 _5468_ (.A(_0802_),
    .B(_2816_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _5469_ (.A(_0804_),
    .B(_0469_),
    .Y(_2175_));
 sky130_fd_sc_hd__nand2_1 _5470_ (.A(_2174_),
    .B(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__a221oi_1 _5471_ (.A1(_2812_),
    .A2(_0800_),
    .B1(_0801_),
    .B2(_0777_),
    .C1(_2176_),
    .Y(_2177_));
 sky130_fd_sc_hd__and4_2 _5472_ (.A(_2167_),
    .B(_2170_),
    .C(_2173_),
    .D(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__nand2_1 _5473_ (.A(_0812_),
    .B(_2907_),
    .Y(_2179_));
 sky130_fd_sc_hd__o21ai_1 _5474_ (.A1(_0337_),
    .A2(_0811_),
    .B1(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__a221oi_1 _5475_ (.A1(_2800_),
    .A2(_0809_),
    .B1(_2814_),
    .B2(_0810_),
    .C1(_2180_),
    .Y(_2181_));
 sky130_fd_sc_hd__nand2_1 _5476_ (.A(_0818_),
    .B(_0886_),
    .Y(_2182_));
 sky130_fd_sc_hd__nand2_1 _5477_ (.A(_0820_),
    .B(_0625_),
    .Y(_2183_));
 sky130_fd_sc_hd__nand2_1 _5478_ (.A(_2182_),
    .B(_2183_),
    .Y(_2184_));
 sky130_fd_sc_hd__a221oi_1 _5479_ (.A1(_0816_),
    .A2(_2806_),
    .B1(_0817_),
    .B2(_2874_),
    .C1(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__o22ai_1 _5480_ (.A1(_3091_),
    .A2(_0826_),
    .B1(_0480_),
    .B2(_0827_),
    .Y(_2186_));
 sky130_fd_sc_hd__a221oi_1 _5481_ (.A1(_0824_),
    .A2(_2935_),
    .B1(_0825_),
    .B2(_0378_),
    .C1(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__nand2_1 _5482_ (.A(_0833_),
    .B(_0458_),
    .Y(_2188_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_0835_),
    .B(_1116_),
    .Y(_2189_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_2188_),
    .B(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__a221oi_1 _5485_ (.A1(_0477_),
    .A2(_0831_),
    .B1(_0832_),
    .B2(_1011_),
    .C1(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__and4_1 _5486_ (.A(_2181_),
    .B(_2185_),
    .C(_2187_),
    .D(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(_0844_),
    .B(_3066_),
    .Y(_2193_));
 sky130_fd_sc_hd__o21ai_1 _5488_ (.A1(_0602_),
    .A2(_0843_),
    .B1(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__a221oi_1 _5489_ (.A1(_3007_),
    .A2(_0840_),
    .B1(_0406_),
    .B2(_0842_),
    .C1(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hd__nand2_1 _5490_ (.A(_2866_),
    .B(_0343_),
    .Y(_2196_));
 sky130_fd_sc_hd__o21ai_1 _5491_ (.A1(_3011_),
    .A2(_0850_),
    .B1(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__a221oi_1 _5492_ (.A1(_2920_),
    .A2(_0848_),
    .B1(_3097_),
    .B2(_0849_),
    .C1(_2197_),
    .Y(_2198_));
 sky130_fd_sc_hd__nand2_1 _5493_ (.A(_2857_),
    .B(_0587_),
    .Y(_2199_));
 sky130_fd_sc_hd__o21ai_1 _5494_ (.A1(_3154_),
    .A2(_2853_),
    .B1(_2199_),
    .Y(_2200_));
 sky130_fd_sc_hd__a221oi_1 _5495_ (.A1(_0742_),
    .A2(_2839_),
    .B1(_2846_),
    .B2(_0871_),
    .C1(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__o22ai_1 _5496_ (.A1(_0349_),
    .A2(_2911_),
    .B1(_3144_),
    .B2(_2916_),
    .Y(_2202_));
 sky130_fd_sc_hd__a221oi_1 _5497_ (.A1(_2974_),
    .A2(_0857_),
    .B1(_0333_),
    .B2(_0858_),
    .C1(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__and4_1 _5498_ (.A(_2195_),
    .B(_2198_),
    .C(_2201_),
    .D(_2203_),
    .X(_2204_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_0865_),
    .B(_0346_),
    .Y(_2205_));
 sky130_fd_sc_hd__nand2_1 _5500_ (.A(_0867_),
    .B(_0392_),
    .Y(_2206_));
 sky130_fd_sc_hd__nand2_1 _5501_ (.A(_2205_),
    .B(_2206_),
    .Y(_2207_));
 sky130_fd_sc_hd__a221oi_2 _5502_ (.A1(_3142_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_2951_),
    .C1(_2207_),
    .Y(_2208_));
 sky130_fd_sc_hd__nand2_1 _5503_ (.A(_0874_),
    .B(_0443_),
    .Y(_2209_));
 sky130_fd_sc_hd__nand2_1 _5504_ (.A(_0877_),
    .B(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .Y(_2210_));
 sky130_fd_sc_hd__nand2_1 _5505_ (.A(_2209_),
    .B(_2210_),
    .Y(_2211_));
 sky130_fd_sc_hd__a221oi_1 _5506_ (.A1(_3002_),
    .A2(_0872_),
    .B1(_0420_),
    .B2(_0873_),
    .C1(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__nand2_1 _5507_ (.A(_0895_),
    .B(_0988_),
    .Y(_2213_));
 sky130_fd_sc_hd__nand2_1 _5508_ (.A(_0897_),
    .B(_0920_),
    .Y(_2214_));
 sky130_fd_sc_hd__nand2_1 _5509_ (.A(_2213_),
    .B(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__a221oi_1 _5510_ (.A1(_0892_),
    .A2(_0894_),
    .B1(_0893_),
    .B2(_0607_),
    .C1(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__nand2_1 _5511_ (.A(_0883_),
    .B(_2887_),
    .Y(_2217_));
 sky130_fd_sc_hd__nand2_1 _5512_ (.A(_0885_),
    .B(_0414_),
    .Y(_2218_));
 sky130_fd_sc_hd__or2b_1 _5513_ (.A(_0889_),
    .B_N(\egd_top.BitStream_buffer.BS_buffer[75] ),
    .X(_2219_));
 sky130_fd_sc_hd__o2111a_1 _5514_ (.A1(_0983_),
    .A2(_0882_),
    .B1(_2217_),
    .C1(_2218_),
    .D1(_2219_),
    .X(_2220_));
 sky130_fd_sc_hd__and4_1 _5515_ (.A(_2208_),
    .B(_2212_),
    .C(_2216_),
    .D(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__and4_1 _5516_ (.A(_2178_),
    .B(_2192_),
    .C(_2204_),
    .D(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__o22ai_1 _5517_ (.A1(_1287_),
    .A2(_0404_),
    .B1(_0641_),
    .B2(_0408_),
    .Y(_2223_));
 sky130_fd_sc_hd__a221oi_1 _5518_ (.A1(_0981_),
    .A2(_2913_),
    .B1(_0982_),
    .B2(_2980_),
    .C1(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__nand2_1 _5519_ (.A(_0990_),
    .B(_2990_),
    .Y(_2225_));
 sky130_fd_sc_hd__nand2_1 _5520_ (.A(_0992_),
    .B(_3070_),
    .Y(_2226_));
 sky130_fd_sc_hd__nand2_1 _5521_ (.A(_2225_),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a221oi_1 _5522_ (.A1(_3015_),
    .A2(_0987_),
    .B1(_2993_),
    .B2(_0989_),
    .C1(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(_0427_),
    .B(\egd_top.BitStream_buffer.BS_buffer[90] ),
    .Y(_2229_));
 sky130_fd_sc_hd__nand2_1 _5524_ (.A(_0999_),
    .B(\egd_top.BitStream_buffer.BS_buffer[94] ),
    .Y(_2230_));
 sky130_fd_sc_hd__nand2_1 _5525_ (.A(_2229_),
    .B(_2230_),
    .Y(_2231_));
 sky130_fd_sc_hd__a221oi_1 _5526_ (.A1(\egd_top.BitStream_buffer.BS_buffer[81] ),
    .A2(_0996_),
    .B1(_0830_),
    .B2(_0997_),
    .C1(_2231_),
    .Y(_2232_));
 sky130_fd_sc_hd__a22o_1 _5527_ (.A1(_0438_),
    .A2(_3037_),
    .B1(_0440_),
    .B2(_3053_),
    .X(_2233_));
 sky130_fd_sc_hd__o22ai_1 _5528_ (.A1(_0957_),
    .A2(_0445_),
    .B1(_1017_),
    .B2(_0448_),
    .Y(_2234_));
 sky130_fd_sc_hd__nor2_1 _5529_ (.A(_2233_),
    .B(_2234_),
    .Y(_2235_));
 sky130_fd_sc_hd__and4_1 _5530_ (.A(_2224_),
    .B(_2228_),
    .C(_2232_),
    .D(_2235_),
    .X(_2236_));
 sky130_fd_sc_hd__nand2_1 _5531_ (.A(_3117_),
    .B(_0366_),
    .Y(_2237_));
 sky130_fd_sc_hd__o21ai_1 _5532_ (.A1(_1533_),
    .A2(_3109_),
    .B1(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__a221oi_1 _5533_ (.A1(_0398_),
    .A2(_0907_),
    .B1(_0553_),
    .B2(_0908_),
    .C1(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__nand2_1 _5534_ (.A(_3099_),
    .B(_0402_),
    .Y(_2240_));
 sky130_fd_sc_hd__o21ai_1 _5535_ (.A1(_3133_),
    .A2(_3092_),
    .B1(_2240_),
    .Y(_2241_));
 sky130_fd_sc_hd__a221oi_2 _5536_ (.A1(_3146_),
    .A2(_3095_),
    .B1(_3103_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[85] ),
    .C1(_2241_),
    .Y(_2242_));
 sky130_fd_sc_hd__or2_1 _5537_ (.A(_0601_),
    .B(_3079_),
    .X(_2243_));
 sky130_fd_sc_hd__or2_1 _5538_ (.A(_0984_),
    .B(_3083_),
    .X(_2244_));
 sky130_fd_sc_hd__nand2_1 _5539_ (.A(_3086_),
    .B(_2957_),
    .Y(_2245_));
 sky130_fd_sc_hd__o2111a_1 _5540_ (.A1(_1301_),
    .A2(_3076_),
    .B1(_2243_),
    .C1(_2244_),
    .D1(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__a22o_1 _5541_ (.A1(_3122_),
    .A2(_2939_),
    .B1(_3125_),
    .B2(_2931_),
    .X(_2247_));
 sky130_fd_sc_hd__o22ai_1 _5542_ (.A1(_1647_),
    .A2(_3130_),
    .B1(_0904_),
    .B2(_3134_),
    .Y(_2248_));
 sky130_fd_sc_hd__nor2_1 _5543_ (.A(_2247_),
    .B(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__and4_1 _5544_ (.A(_2239_),
    .B(_2242_),
    .C(_2246_),
    .D(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__and2_1 _5545_ (.A(_2236_),
    .B(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__a22o_1 _5546_ (.A1(_0495_),
    .A2(_0930_),
    .B1(_0931_),
    .B2(_1000_),
    .X(_2252_));
 sky130_fd_sc_hd__a221oi_1 _5547_ (.A1(_3034_),
    .A2(_0933_),
    .B1(_3048_),
    .B2(_0934_),
    .C1(_2252_),
    .Y(_2253_));
 sky130_fd_sc_hd__nand2_1 _5548_ (.A(_0925_),
    .B(_0638_),
    .Y(_2254_));
 sky130_fd_sc_hd__o21ai_1 _5549_ (.A1(_0619_),
    .A2(_0923_),
    .B1(_2254_),
    .Y(_2255_));
 sky130_fd_sc_hd__a221oi_2 _5550_ (.A1(_0610_),
    .A2(_0921_),
    .B1(_3030_),
    .B2(_0922_),
    .C1(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__nand2_1 _5551_ (.A(_0939_),
    .B(_2926_),
    .Y(_2257_));
 sky130_fd_sc_hd__nand2_1 _5552_ (.A(_0941_),
    .B(_2959_),
    .Y(_2258_));
 sky130_fd_sc_hd__nand2_1 _5553_ (.A(_2257_),
    .B(_2258_),
    .Y(_2259_));
 sky130_fd_sc_hd__a221oi_1 _5554_ (.A1(_0937_),
    .A2(_2859_),
    .B1(_0463_),
    .B2(_0938_),
    .C1(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__nand2_1 _5555_ (.A(_0947_),
    .B(_3105_),
    .Y(_2261_));
 sky130_fd_sc_hd__nand2_1 _5556_ (.A(_0949_),
    .B(_0709_),
    .Y(_2262_));
 sky130_fd_sc_hd__nand2_1 _5557_ (.A(_2261_),
    .B(_2262_),
    .Y(_2263_));
 sky130_fd_sc_hd__a221oi_1 _5558_ (.A1(_0875_),
    .A2(_0945_),
    .B1(_0946_),
    .B2(_3112_),
    .C1(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__and4_1 _5559_ (.A(_2253_),
    .B(_2256_),
    .C(_2260_),
    .D(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__o22ai_2 _5560_ (.A1(_0723_),
    .A2(_0956_),
    .B1(_1717_),
    .B2(_0958_),
    .Y(_2266_));
 sky130_fd_sc_hd__a221oi_4 _5561_ (.A1(_2826_),
    .A2(_0954_),
    .B1(_2824_),
    .B2(_0955_),
    .C1(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__o22ai_1 _5562_ (.A1(_3129_),
    .A2(_0963_),
    .B1(_0717_),
    .B2(_0964_),
    .Y(_2268_));
 sky130_fd_sc_hd__a221oi_1 _5563_ (.A1(_0464_),
    .A2(_0961_),
    .B1(_0962_),
    .B2(_2848_),
    .C1(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__o22ai_1 _5564_ (.A1(_0888_),
    .A2(_0969_),
    .B1(_1075_),
    .B2(_0971_),
    .Y(_2270_));
 sky130_fd_sc_hd__a221oi_1 _5565_ (.A1(_0967_),
    .A2(_2881_),
    .B1(_0968_),
    .B2(_2943_),
    .C1(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__o22ai_1 _5566_ (.A1(_3108_),
    .A2(_0976_),
    .B1(_0561_),
    .B2(_0977_),
    .Y(_2272_));
 sky130_fd_sc_hd__a221oi_1 _5567_ (.A1(_0974_),
    .A2(_3119_),
    .B1(_0975_),
    .B2(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .C1(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__and4_1 _5568_ (.A(_2267_),
    .B(_2269_),
    .C(_2271_),
    .D(_2273_),
    .X(_2274_));
 sky130_fd_sc_hd__and3_1 _5569_ (.A(_2251_),
    .B(_2265_),
    .C(_2274_),
    .X(_2275_));
 sky130_fd_sc_hd__nand3_2 _5570_ (.A(_2222_),
    .B(_0903_),
    .C(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__o21a_1 _5571_ (.A1(_0412_),
    .A2(_0456_),
    .B1(_2789_),
    .X(_2277_));
 sky130_fd_sc_hd__nand2_1 _5572_ (.A(_2276_),
    .B(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__nand2_1 _5573_ (.A(net221),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2279_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(_2278_),
    .B(_2279_),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_2 _5575_ (.A(_2793_),
    .B(_2776_),
    .Y(_2280_));
 sky130_fd_sc_hd__buf_4 _5576_ (.A(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__mux2_1 _5577_ (.A0(net7),
    .A1(_0458_),
    .S(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__clkbuf_1 _5578_ (.A(_2282_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _5579_ (.A0(net6),
    .A1(_0625_),
    .S(_2281_),
    .X(_2283_));
 sky130_fd_sc_hd__clkbuf_1 _5580_ (.A(_2283_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _5581_ (.A0(net5),
    .A1(_0777_),
    .S(_2281_),
    .X(_2284_));
 sky130_fd_sc_hd__clkbuf_1 _5582_ (.A(_2284_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(net4),
    .A1(_1011_),
    .S(_2281_),
    .X(_2285_));
 sky130_fd_sc_hd__clkbuf_1 _5584_ (.A(_2285_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _5585_ (.A0(net3),
    .A1(_0886_),
    .S(_2281_),
    .X(_2286_));
 sky130_fd_sc_hd__clkbuf_1 _5586_ (.A(_2286_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(net2),
    .A1(_2874_),
    .S(_2281_),
    .X(_2287_));
 sky130_fd_sc_hd__clkbuf_1 _5588_ (.A(_2287_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(net16),
    .A1(_0469_),
    .S(_2281_),
    .X(_2288_));
 sky130_fd_sc_hd__clkbuf_1 _5590_ (.A(_2288_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(net15),
    .A1(_0988_),
    .S(_2281_),
    .X(_2289_));
 sky130_fd_sc_hd__clkbuf_1 _5592_ (.A(_2289_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(net14),
    .A1(_1116_),
    .S(_2281_),
    .X(_2290_));
 sky130_fd_sc_hd__clkbuf_1 _5594_ (.A(_2290_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5595_ (.A0(net13),
    .A1(_0841_),
    .S(_2281_),
    .X(_2291_));
 sky130_fd_sc_hd__clkbuf_1 _5596_ (.A(_2291_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(net12),
    .A1(_3101_),
    .S(_2281_),
    .X(_2292_));
 sky130_fd_sc_hd__clkbuf_1 _5598_ (.A(_2292_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(net11),
    .A1(_0551_),
    .S(_2281_),
    .X(_2293_));
 sky130_fd_sc_hd__clkbuf_1 _5600_ (.A(_2293_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(net10),
    .A1(_2881_),
    .S(_2280_),
    .X(_2294_));
 sky130_fd_sc_hd__clkbuf_1 _5602_ (.A(_2294_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5603_ (.A0(net9),
    .A1(_2943_),
    .S(_2280_),
    .X(_2295_));
 sky130_fd_sc_hd__clkbuf_1 _5604_ (.A(_2295_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5605_ (.A0(net8),
    .A1(_0412_),
    .S(_2280_),
    .X(_2296_));
 sky130_fd_sc_hd__clkbuf_1 _5606_ (.A(_2296_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5607_ (.A0(net1),
    .A1(_0414_),
    .S(_2280_),
    .X(_2297_));
 sky130_fd_sc_hd__clkbuf_1 _5608_ (.A(_2297_),
    .X(_0274_));
 sky130_fd_sc_hd__or4b_4 _5609_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(_2775_),
    .D_N(_2793_),
    .X(_2298_));
 sky130_fd_sc_hd__buf_4 _5610_ (.A(_2298_),
    .X(_2299_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(net7),
    .A1(_2887_),
    .S(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__clkbuf_1 _5612_ (.A(_2300_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5613_ (.A0(net6),
    .A1(_3007_),
    .S(_2299_),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _5614_ (.A(_2301_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5615_ (.A0(net5),
    .A1(_2993_),
    .S(_2299_),
    .X(_2302_));
 sky130_fd_sc_hd__clkbuf_1 _5616_ (.A(_2302_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5617_ (.A0(net4),
    .A1(_3010_),
    .S(_2299_),
    .X(_2303_));
 sky130_fd_sc_hd__clkbuf_1 _5618_ (.A(_2303_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5619_ (.A0(net3),
    .A1(_0406_),
    .S(_2299_),
    .X(_2304_));
 sky130_fd_sc_hd__clkbuf_1 _5620_ (.A(_2304_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5621_ (.A0(net2),
    .A1(_3040_),
    .S(_2299_),
    .X(_2305_));
 sky130_fd_sc_hd__clkbuf_1 _5622_ (.A(_2305_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5623_ (.A0(net16),
    .A1(_3015_),
    .S(_2299_),
    .X(_2306_));
 sky130_fd_sc_hd__clkbuf_1 _5624_ (.A(_2306_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5625_ (.A0(net15),
    .A1(_3017_),
    .S(_2299_),
    .X(_2307_));
 sky130_fd_sc_hd__clkbuf_1 _5626_ (.A(_2307_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5627_ (.A0(net14),
    .A1(_0402_),
    .S(_2299_),
    .X(_2308_));
 sky130_fd_sc_hd__clkbuf_1 _5628_ (.A(_2308_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5629_ (.A0(net13),
    .A1(_2863_),
    .S(_2299_),
    .X(_2309_));
 sky130_fd_sc_hd__clkbuf_1 _5630_ (.A(_2309_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5631_ (.A0(net12),
    .A1(_2920_),
    .S(_2299_),
    .X(_2310_));
 sky130_fd_sc_hd__clkbuf_1 _5632_ (.A(_2310_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5633_ (.A0(net11),
    .A1(_2922_),
    .S(_2299_),
    .X(_2311_));
 sky130_fd_sc_hd__clkbuf_1 _5634_ (.A(_2311_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5635_ (.A0(net10),
    .A1(_2913_),
    .S(_2298_),
    .X(_2312_));
 sky130_fd_sc_hd__clkbuf_1 _5636_ (.A(_2312_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5637_ (.A0(net9),
    .A1(_2980_),
    .S(_2298_),
    .X(_2313_));
 sky130_fd_sc_hd__clkbuf_1 _5638_ (.A(_2313_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5639_ (.A0(net8),
    .A1(_3097_),
    .S(_2298_),
    .X(_2314_));
 sky130_fd_sc_hd__clkbuf_1 _5640_ (.A(_2314_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5641_ (.A0(net1),
    .A1(_3090_),
    .S(_2298_),
    .X(_2315_));
 sky130_fd_sc_hd__clkbuf_1 _5642_ (.A(_2315_),
    .X(_0258_));
 sky130_fd_sc_hd__or4b_4 _5643_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(_2774_),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .D_N(_2793_),
    .X(_2316_));
 sky130_fd_sc_hd__clkbuf_8 _5644_ (.A(_2316_),
    .X(_2317_));
 sky130_fd_sc_hd__mux2_1 _5645_ (.A0(net7),
    .A1(_2907_),
    .S(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__clkbuf_1 _5646_ (.A(_2318_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5647_ (.A0(net6),
    .A1(_3127_),
    .S(_2317_),
    .X(_2319_));
 sky130_fd_sc_hd__clkbuf_1 _5648_ (.A(_2319_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5649_ (.A0(net5),
    .A1(_3124_),
    .S(_2317_),
    .X(_2320_));
 sky130_fd_sc_hd__clkbuf_1 _5650_ (.A(_2320_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5651_ (.A0(net4),
    .A1(_0395_),
    .S(_2317_),
    .X(_2321_));
 sky130_fd_sc_hd__clkbuf_1 _5652_ (.A(_2321_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5653_ (.A0(net3),
    .A1(_2935_),
    .S(_2317_),
    .X(_2322_));
 sky130_fd_sc_hd__clkbuf_1 _5654_ (.A(_2322_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5655_ (.A0(net2),
    .A1(_0378_),
    .S(_2317_),
    .X(_2323_));
 sky130_fd_sc_hd__clkbuf_1 _5656_ (.A(_2323_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5657_ (.A0(net16),
    .A1(_0341_),
    .S(_2317_),
    .X(_2324_));
 sky130_fd_sc_hd__clkbuf_1 _5658_ (.A(_2324_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5659_ (.A0(net15),
    .A1(_0343_),
    .S(_2317_),
    .X(_2325_));
 sky130_fd_sc_hd__clkbuf_1 _5660_ (.A(_2325_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5661_ (.A0(net14),
    .A1(_2974_),
    .S(_2317_),
    .X(_2326_));
 sky130_fd_sc_hd__clkbuf_1 _5662_ (.A(_2326_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(net13),
    .A1(_0333_),
    .S(_2317_),
    .X(_2327_));
 sky130_fd_sc_hd__clkbuf_1 _5664_ (.A(_2327_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5665_ (.A0(net12),
    .A1(_3143_),
    .S(_2317_),
    .X(_2328_));
 sky130_fd_sc_hd__clkbuf_1 _5666_ (.A(_2328_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5667_ (.A0(net11),
    .A1(_0336_),
    .S(_2317_),
    .X(_2329_));
 sky130_fd_sc_hd__clkbuf_1 _5668_ (.A(_2329_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(net10),
    .A1(_3146_),
    .S(_2316_),
    .X(_2330_));
 sky130_fd_sc_hd__clkbuf_1 _5670_ (.A(_2330_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5671_ (.A0(net9),
    .A1(_3132_),
    .S(_2316_),
    .X(_2331_));
 sky130_fd_sc_hd__clkbuf_1 _5672_ (.A(_2331_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5673_ (.A0(net8),
    .A1(\egd_top.BitStream_buffer.BS_buffer[46] ),
    .S(_2316_),
    .X(_2332_));
 sky130_fd_sc_hd__clkbuf_1 _5674_ (.A(_2332_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5675_ (.A0(net1),
    .A1(_2931_),
    .S(_2316_),
    .X(_2333_));
 sky130_fd_sc_hd__clkbuf_1 _5676_ (.A(_2333_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_4 _5677_ (.A(\egd_top.BitStream_buffer.buffer_index[6] ),
    .B(_2795_),
    .X(_2334_));
 sky130_fd_sc_hd__buf_4 _5678_ (.A(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__mux2_1 _5679_ (.A0(net7),
    .A1(_2939_),
    .S(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__clkbuf_1 _5680_ (.A(_2336_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5681_ (.A0(net6),
    .A1(_2926_),
    .S(_2335_),
    .X(_2337_));
 sky130_fd_sc_hd__clkbuf_1 _5682_ (.A(_2337_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5683_ (.A0(net5),
    .A1(_0346_),
    .S(_2335_),
    .X(_2338_));
 sky130_fd_sc_hd__clkbuf_1 _5684_ (.A(_2338_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5685_ (.A0(net4),
    .A1(_3112_),
    .S(_2335_),
    .X(_2339_));
 sky130_fd_sc_hd__clkbuf_1 _5686_ (.A(_2339_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _5687_ (.A0(net3),
    .A1(_3119_),
    .S(_2335_),
    .X(_2340_));
 sky130_fd_sc_hd__clkbuf_1 _5688_ (.A(_2340_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5689_ (.A0(net2),
    .A1(\egd_top.BitStream_buffer.BS_buffer[53] ),
    .S(_2335_),
    .X(_2341_));
 sky130_fd_sc_hd__clkbuf_1 _5690_ (.A(_2341_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(net16),
    .A1(\egd_top.BitStream_buffer.BS_buffer[54] ),
    .S(_2335_),
    .X(_2342_));
 sky130_fd_sc_hd__clkbuf_1 _5692_ (.A(_2342_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5693_ (.A0(net15),
    .A1(\egd_top.BitStream_buffer.BS_buffer[55] ),
    .S(_2335_),
    .X(_2343_));
 sky130_fd_sc_hd__clkbuf_1 _5694_ (.A(_2343_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5695_ (.A0(net14),
    .A1(\egd_top.BitStream_buffer.BS_buffer[56] ),
    .S(_2335_),
    .X(_2344_));
 sky130_fd_sc_hd__clkbuf_1 _5696_ (.A(_2344_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(net13),
    .A1(\egd_top.BitStream_buffer.BS_buffer[57] ),
    .S(_2335_),
    .X(_2345_));
 sky130_fd_sc_hd__clkbuf_1 _5698_ (.A(_2345_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5699_ (.A0(net12),
    .A1(_3115_),
    .S(_2335_),
    .X(_2346_));
 sky130_fd_sc_hd__clkbuf_1 _5700_ (.A(_2346_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5701_ (.A0(net11),
    .A1(_0385_),
    .S(_2335_),
    .X(_2347_));
 sky130_fd_sc_hd__clkbuf_1 _5702_ (.A(_2347_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5703_ (.A0(net10),
    .A1(_0389_),
    .S(_2334_),
    .X(_2348_));
 sky130_fd_sc_hd__clkbuf_1 _5704_ (.A(_2348_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(net9),
    .A1(_2951_),
    .S(_2334_),
    .X(_2349_));
 sky130_fd_sc_hd__clkbuf_1 _5706_ (.A(_2349_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(net8),
    .A1(_0392_),
    .S(_2334_),
    .X(_2350_));
 sky130_fd_sc_hd__clkbuf_1 _5708_ (.A(_2350_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(net1),
    .A1(_3142_),
    .S(_2334_),
    .X(_2351_));
 sky130_fd_sc_hd__clkbuf_1 _5710_ (.A(_2351_),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_2 _5711_ (.A(_2793_),
    .B(_2779_),
    .Y(_2352_));
 sky130_fd_sc_hd__buf_4 _5712_ (.A(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _5713_ (.A0(net7),
    .A1(_3139_),
    .S(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__clkbuf_1 _5714_ (.A(_2354_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5715_ (.A0(net6),
    .A1(_0398_),
    .S(_2353_),
    .X(_2355_));
 sky130_fd_sc_hd__clkbuf_1 _5716_ (.A(_2355_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5717_ (.A0(net5),
    .A1(_0366_),
    .S(_2353_),
    .X(_2356_));
 sky130_fd_sc_hd__clkbuf_1 _5718_ (.A(_2356_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(net4),
    .A1(_0435_),
    .S(_2353_),
    .X(_2357_));
 sky130_fd_sc_hd__clkbuf_1 _5720_ (.A(_2357_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5721_ (.A0(net3),
    .A1(_2957_),
    .S(_2353_),
    .X(_2358_));
 sky130_fd_sc_hd__clkbuf_1 _5722_ (.A(_2358_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5723_ (.A0(net2),
    .A1(_0371_),
    .S(_2353_),
    .X(_2359_));
 sky130_fd_sc_hd__clkbuf_1 _5724_ (.A(_2359_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5725_ (.A0(net16),
    .A1(_0656_),
    .S(_2353_),
    .X(_2360_));
 sky130_fd_sc_hd__clkbuf_1 _5726_ (.A(_2360_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(net15),
    .A1(_3105_),
    .S(_2353_),
    .X(_2361_));
 sky130_fd_sc_hd__clkbuf_1 _5728_ (.A(_2361_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(net14),
    .A1(_0553_),
    .S(_2353_),
    .X(_2362_));
 sky130_fd_sc_hd__clkbuf_1 _5730_ (.A(_2362_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _5731_ (.A0(net13),
    .A1(_0709_),
    .S(_2353_),
    .X(_2363_));
 sky130_fd_sc_hd__clkbuf_1 _5732_ (.A(_2363_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5733_ (.A0(net12),
    .A1(_2859_),
    .S(_2353_),
    .X(_2364_));
 sky130_fd_sc_hd__clkbuf_1 _5734_ (.A(_2364_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5735_ (.A0(net11),
    .A1(_2830_),
    .S(_2353_),
    .X(_2365_));
 sky130_fd_sc_hd__clkbuf_1 _5736_ (.A(_2365_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _5737_ (.A0(net10),
    .A1(_0463_),
    .S(_2352_),
    .X(_2366_));
 sky130_fd_sc_hd__clkbuf_1 _5738_ (.A(_2366_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5739_ (.A0(net9),
    .A1(_2848_),
    .S(_2352_),
    .X(_2367_));
 sky130_fd_sc_hd__clkbuf_1 _5740_ (.A(_2367_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(net8),
    .A1(_0464_),
    .S(_2352_),
    .X(_2368_));
 sky130_fd_sc_hd__clkbuf_1 _5742_ (.A(_2368_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _5743_ (.A0(net1),
    .A1(_2959_),
    .S(_2352_),
    .X(_2369_));
 sky130_fd_sc_hd__clkbuf_1 _5744_ (.A(_2369_),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _5745_ (.A(_2795_),
    .B(_2773_),
    .Y(_2370_));
 sky130_fd_sc_hd__and2_1 _5746_ (.A(_2798_),
    .B(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__clkbuf_1 _5747_ (.A(_2371_),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(_2794_),
    .B(_2774_),
    .Y(_2372_));
 sky130_fd_sc_hd__and2_1 _5749_ (.A(_2795_),
    .B(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__clkbuf_1 _5750_ (.A(_2373_),
    .X(_0208_));
 sky130_fd_sc_hd__or2_1 _5751_ (.A(\egd_top.BitStream_buffer.buffer_index[4] ),
    .B(net224),
    .X(_2374_));
 sky130_fd_sc_hd__and2_1 _5752_ (.A(_2374_),
    .B(_2794_),
    .X(_2375_));
 sky130_fd_sc_hd__clkbuf_1 _5753_ (.A(_2375_),
    .X(_0207_));
 sky130_fd_sc_hd__or4b_4 _5754_ (.A(_2773_),
    .B(_2774_),
    .C(\egd_top.BitStream_buffer.buffer_index[4] ),
    .D_N(_2793_),
    .X(_2376_));
 sky130_fd_sc_hd__buf_4 _5755_ (.A(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_1 _5756_ (.A0(net7),
    .A1(_0638_),
    .S(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__clkbuf_1 _5757_ (.A(_2378_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(net6),
    .A1(_0610_),
    .S(_2377_),
    .X(_2379_));
 sky130_fd_sc_hd__clkbuf_1 _5759_ (.A(_2379_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _5760_ (.A0(net5),
    .A1(_0443_),
    .S(_2377_),
    .X(_2380_));
 sky130_fd_sc_hd__clkbuf_1 _5761_ (.A(_2380_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(net4),
    .A1(_2987_),
    .S(_2377_),
    .X(_2381_));
 sky130_fd_sc_hd__clkbuf_1 _5763_ (.A(_2381_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(net3),
    .A1(_3034_),
    .S(_2377_),
    .X(_2382_));
 sky130_fd_sc_hd__clkbuf_1 _5765_ (.A(_2382_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(net2),
    .A1(_3048_),
    .S(_2377_),
    .X(_2383_));
 sky130_fd_sc_hd__clkbuf_1 _5767_ (.A(_2383_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(net16),
    .A1(_3002_),
    .S(_2377_),
    .X(_2384_));
 sky130_fd_sc_hd__clkbuf_1 _5769_ (.A(_2384_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _5770_ (.A0(net15),
    .A1(_3030_),
    .S(_2377_),
    .X(_2385_));
 sky130_fd_sc_hd__clkbuf_1 _5771_ (.A(_2385_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(net14),
    .A1(_3037_),
    .S(_2377_),
    .X(_2386_));
 sky130_fd_sc_hd__clkbuf_1 _5773_ (.A(_2386_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(net13),
    .A1(_3053_),
    .S(_2377_),
    .X(_2387_));
 sky130_fd_sc_hd__clkbuf_1 _5775_ (.A(_2387_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5776_ (.A0(net12),
    .A1(_2990_),
    .S(_2377_),
    .X(_2388_));
 sky130_fd_sc_hd__clkbuf_1 _5777_ (.A(_2388_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _5778_ (.A0(net11),
    .A1(_3058_),
    .S(_2377_),
    .X(_2389_));
 sky130_fd_sc_hd__clkbuf_1 _5779_ (.A(_2389_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _5780_ (.A0(net10),
    .A1(_3066_),
    .S(_2376_),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_1 _5781_ (.A(_2390_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(net9),
    .A1(_3153_),
    .S(_2376_),
    .X(_2391_));
 sky130_fd_sc_hd__clkbuf_1 _5783_ (.A(_2391_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(net8),
    .A1(_3070_),
    .S(_2376_),
    .X(_2392_));
 sky130_fd_sc_hd__clkbuf_1 _5785_ (.A(_2392_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _5786_ (.A0(net1),
    .A1(_0330_),
    .S(_2376_),
    .X(_2393_));
 sky130_fd_sc_hd__clkbuf_1 _5787_ (.A(_2393_),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _5788_ (.A(\egd_top.BitStream_buffer.pc_reg[5] ),
    .Y(_2394_));
 sky130_fd_sc_hd__or2_1 _5789_ (.A(\egd_top.BitStream_buffer.pc_reg[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .X(_2395_));
 sky130_fd_sc_hd__nand2_1 _5790_ (.A(\egd_top.BitStream_buffer.pc_reg[1] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[1] ),
    .Y(_2396_));
 sky130_fd_sc_hd__nand2_2 _5791_ (.A(_2395_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__o21ai_4 _5792_ (.A1(_2762_),
    .A2(_2397_),
    .B1(_2396_),
    .Y(_2398_));
 sky130_fd_sc_hd__or2_1 _5793_ (.A(\egd_top.BitStream_buffer.pc_reg[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .X(_2399_));
 sky130_fd_sc_hd__nand2_1 _5794_ (.A(\egd_top.BitStream_buffer.pc_reg[2] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[2] ),
    .Y(_2400_));
 sky130_fd_sc_hd__a21bo_2 _5795_ (.A1(_2398_),
    .A2(_2399_),
    .B1_N(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__or2_1 _5796_ (.A(\egd_top.BitStream_buffer.pc_reg[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .X(_2402_));
 sky130_fd_sc_hd__nand2_1 _5797_ (.A(\egd_top.BitStream_buffer.pc_reg[3] ),
    .B(\egd_top.BitStream_buffer.exp_golomb_len[3] ),
    .Y(_2403_));
 sky130_fd_sc_hd__a21bo_1 _5798_ (.A1(_2401_),
    .A2(_2402_),
    .B1_N(_2403_),
    .X(_2404_));
 sky130_fd_sc_hd__nand2_1 _5799_ (.A(_2404_),
    .B(\egd_top.BitStream_buffer.pc_reg[4] ),
    .Y(_2405_));
 sky130_fd_sc_hd__nor2_2 _5800_ (.A(_2394_),
    .B(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__xor2_4 _5801_ (.A(\egd_top.BitStream_buffer.pc_reg[6] ),
    .B(_2406_),
    .X(\egd_top.BitStream_buffer.pc[6] ));
 sky130_fd_sc_hd__nand2_1 _5802_ (.A(net35),
    .B(\egd_top.BitStream_buffer.pc[6] ),
    .Y(_2407_));
 sky130_fd_sc_hd__inv_2 _5803_ (.A(_2407_),
    .Y(_0190_));
 sky130_fd_sc_hd__and2_1 _5804_ (.A(_2405_),
    .B(_2394_),
    .X(_2408_));
 sky130_fd_sc_hd__nor2_2 _5805_ (.A(_2406_),
    .B(_2408_),
    .Y(\egd_top.BitStream_buffer.pc[5] ));
 sky130_fd_sc_hd__nand2_1 _5806_ (.A(net36),
    .B(\egd_top.BitStream_buffer.pc[5] ),
    .Y(_2409_));
 sky130_fd_sc_hd__inv_2 _5807_ (.A(_2409_),
    .Y(_0189_));
 sky130_fd_sc_hd__or2_1 _5808_ (.A(\egd_top.BitStream_buffer.pc_reg[4] ),
    .B(_2404_),
    .X(_2410_));
 sky130_fd_sc_hd__and2_1 _5809_ (.A(_2410_),
    .B(_2405_),
    .X(_2411_));
 sky130_fd_sc_hd__buf_2 _5810_ (.A(_2411_),
    .X(\egd_top.BitStream_buffer.pc[4] ));
 sky130_fd_sc_hd__nand2_1 _5811_ (.A(net36),
    .B(\egd_top.BitStream_buffer.pc[4] ),
    .Y(_2412_));
 sky130_fd_sc_hd__inv_2 _5812_ (.A(_2412_),
    .Y(_0188_));
 sky130_fd_sc_hd__nand2_2 _5813_ (.A(_2402_),
    .B(_2403_),
    .Y(_2413_));
 sky130_fd_sc_hd__xnor2_4 _5814_ (.A(_2413_),
    .B(_2401_),
    .Y(\egd_top.BitStream_buffer.pc[3] ));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(net36),
    .B(\egd_top.BitStream_buffer.pc[3] ),
    .Y(_2414_));
 sky130_fd_sc_hd__inv_2 _5816_ (.A(_2414_),
    .Y(_0187_));
 sky130_fd_sc_hd__nand2_2 _5817_ (.A(_2399_),
    .B(_2400_),
    .Y(_2415_));
 sky130_fd_sc_hd__xnor2_4 _5818_ (.A(_2415_),
    .B(_2398_),
    .Y(\egd_top.BitStream_buffer.pc[2] ));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(net35),
    .B(\egd_top.BitStream_buffer.pc[2] ),
    .Y(_2416_));
 sky130_fd_sc_hd__inv_2 _5820_ (.A(_2416_),
    .Y(_0186_));
 sky130_fd_sc_hd__xor2_4 _5821_ (.A(_2762_),
    .B(_2397_),
    .X(\egd_top.BitStream_buffer.pc[1] ));
 sky130_fd_sc_hd__nand2_1 _5822_ (.A(net37),
    .B(\egd_top.BitStream_buffer.pc[1] ),
    .Y(_2417_));
 sky130_fd_sc_hd__inv_2 _5823_ (.A(_2417_),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(\egd_top.BitStream_buffer.pc[0] ),
    .B(net38),
    .Y(_2418_));
 sky130_fd_sc_hd__inv_2 _5825_ (.A(_2418_),
    .Y(_0184_));
 sky130_fd_sc_hd__or4b_4 _5826_ (.A(_2773_),
    .B(\egd_top.BitStream_buffer.buffer_index[5] ),
    .C(_2775_),
    .D_N(_2793_),
    .X(_2419_));
 sky130_fd_sc_hd__buf_4 _5827_ (.A(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(net7),
    .A1(_0495_),
    .S(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__clkbuf_1 _5829_ (.A(_2421_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _5830_ (.A0(net6),
    .A1(_0657_),
    .S(_2420_),
    .X(_2422_));
 sky130_fd_sc_hd__clkbuf_1 _5831_ (.A(_2422_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(net5),
    .A1(_0894_),
    .S(_2420_),
    .X(_2423_));
 sky130_fd_sc_hd__clkbuf_1 _5833_ (.A(_2423_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _5834_ (.A0(net4),
    .A1(_1000_),
    .S(_2420_),
    .X(_2424_));
 sky130_fd_sc_hd__clkbuf_1 _5835_ (.A(_2424_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(net3),
    .A1(_0830_),
    .S(_2420_),
    .X(_2425_));
 sky130_fd_sc_hd__clkbuf_1 _5837_ (.A(_2425_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _5838_ (.A0(net2),
    .A1(_0926_),
    .S(_2420_),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _5839_ (.A(_2426_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _5840_ (.A0(net16),
    .A1(_0920_),
    .S(_2420_),
    .X(_2427_));
 sky130_fd_sc_hd__clkbuf_1 _5841_ (.A(_2427_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _5842_ (.A0(net15),
    .A1(_0875_),
    .S(_2420_),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_1 _5843_ (.A(_2428_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(net14),
    .A1(_0587_),
    .S(_2420_),
    .X(_2429_));
 sky130_fd_sc_hd__clkbuf_1 _5845_ (.A(_2429_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _5846_ (.A0(net13),
    .A1(_0742_),
    .S(_2420_),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_1 _5847_ (.A(_2430_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5848_ (.A0(net12),
    .A1(_0583_),
    .S(_2420_),
    .X(_2431_));
 sky130_fd_sc_hd__clkbuf_1 _5849_ (.A(_2431_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _5850_ (.A0(net11),
    .A1(_0871_),
    .S(_2420_),
    .X(_2432_));
 sky130_fd_sc_hd__clkbuf_1 _5851_ (.A(_2432_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(net10),
    .A1(_0420_),
    .S(_2419_),
    .X(_2433_));
 sky130_fd_sc_hd__clkbuf_1 _5853_ (.A(_2433_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5854_ (.A0(net9),
    .A1(_0607_),
    .S(_2419_),
    .X(_2434_));
 sky130_fd_sc_hd__clkbuf_1 _5855_ (.A(_2434_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5856_ (.A0(net8),
    .A1(_2904_),
    .S(_2419_),
    .X(_2435_));
 sky130_fd_sc_hd__clkbuf_1 _5857_ (.A(_2435_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(net1),
    .A1(_0477_),
    .S(_2419_),
    .X(_2436_));
 sky130_fd_sc_hd__clkbuf_1 _5859_ (.A(_2436_),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _5860_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2437_));
 sky130_fd_sc_hd__nand2_1 _5861_ (.A(_2437_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2438_));
 sky130_fd_sc_hd__inv_2 _5862_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2439_));
 sky130_fd_sc_hd__nand2_1 _5863_ (.A(_2438_),
    .B(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__inv_2 _5864_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2441_));
 sky130_fd_sc_hd__nand2_1 _5865_ (.A(_2440_),
    .B(_2441_),
    .Y(_2442_));
 sky130_fd_sc_hd__inv_2 _5866_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2443_));
 sky130_fd_sc_hd__nand2_1 _5867_ (.A(_2442_),
    .B(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__inv_2 _5868_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2445_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(_2444_),
    .B(_2445_),
    .Y(_2446_));
 sky130_fd_sc_hd__inv_2 _5870_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2447_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(_2446_),
    .B(_2447_),
    .Y(_2448_));
 sky130_fd_sc_hd__inv_2 _5872_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_2449_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(_2448_),
    .B(_2449_),
    .Y(_2450_));
 sky130_fd_sc_hd__inv_2 _5874_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2451_));
 sky130_fd_sc_hd__nand2_1 _5875_ (.A(_2450_),
    .B(_2451_),
    .Y(_2452_));
 sky130_fd_sc_hd__inv_2 _5876_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2453_));
 sky130_fd_sc_hd__inv_4 _5877_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .Y(_2454_));
 sky130_fd_sc_hd__nand2_1 _5878_ (.A(_2453_),
    .B(_2454_),
    .Y(_2455_));
 sky130_fd_sc_hd__nor2_1 _5879_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hd__inv_2 _5880_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .Y(_2457_));
 sky130_fd_sc_hd__nand2_1 _5881_ (.A(_2456_),
    .B(_2457_),
    .Y(_2458_));
 sky130_fd_sc_hd__inv_2 _5882_ (.A(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__nand2_1 _5883_ (.A(_2452_),
    .B(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__a21oi_1 _5884_ (.A1(_2453_),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2461_));
 sky130_fd_sc_hd__nand2_1 _5885_ (.A(_2460_),
    .B(_2461_),
    .Y(_2462_));
 sky130_fd_sc_hd__nor2_1 _5886_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .Y(_2463_));
 sky130_fd_sc_hd__nand2_1 _5887_ (.A(_2462_),
    .B(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__nor2_1 _5888_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ),
    .Y(_2465_));
 sky130_fd_sc_hd__nand2_2 _5889_ (.A(_2464_),
    .B(_2465_),
    .Y(_2466_));
 sky130_fd_sc_hd__nor2_1 _5890_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2467_));
 sky130_fd_sc_hd__inv_2 _5891_ (.A(_2467_),
    .Y(_2468_));
 sky130_fd_sc_hd__nor2_1 _5892_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B(_2468_),
    .Y(_2469_));
 sky130_fd_sc_hd__inv_2 _5893_ (.A(_2469_),
    .Y(_2470_));
 sky130_fd_sc_hd__and3_1 _5894_ (.A(_2459_),
    .B(_2451_),
    .C(_2449_),
    .X(_2471_));
 sky130_fd_sc_hd__o21ai_1 _5895_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .A2(_2470_),
    .B1(_2471_),
    .Y(_2472_));
 sky130_fd_sc_hd__nand2_1 _5896_ (.A(_2463_),
    .B(_2789_),
    .Y(_2473_));
 sky130_fd_sc_hd__inv_2 _5897_ (.A(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__nor2_1 _5898_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .Y(_2475_));
 sky130_fd_sc_hd__nand2_1 _5899_ (.A(_2474_),
    .B(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__inv_2 _5900_ (.A(_2476_),
    .Y(_2477_));
 sky130_fd_sc_hd__nand2_1 _5901_ (.A(_2472_),
    .B(_2477_),
    .Y(_2478_));
 sky130_fd_sc_hd__inv_2 _5902_ (.A(_2478_),
    .Y(_2479_));
 sky130_fd_sc_hd__nand2_2 _5903_ (.A(_2471_),
    .B(_2474_),
    .Y(_2480_));
 sky130_fd_sc_hd__nand2_4 _5904_ (.A(_2479_),
    .B(_2480_),
    .Y(_2481_));
 sky130_fd_sc_hd__inv_2 _5905_ (.A(_2481_),
    .Y(_2482_));
 sky130_fd_sc_hd__o21a_1 _5906_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .A2(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .B1(_2441_),
    .X(_2483_));
 sky130_fd_sc_hd__a211o_1 _5907_ (.A1(_2483_),
    .A2(_2443_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .C1(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .X(_2484_));
 sky130_fd_sc_hd__nand2_1 _5908_ (.A(_2484_),
    .B(_2471_),
    .Y(_2485_));
 sky130_fd_sc_hd__a21o_1 _5909_ (.A1(_2458_),
    .A2(_2475_),
    .B1(_2473_),
    .X(_2486_));
 sky130_fd_sc_hd__inv_2 _5910_ (.A(_2486_),
    .Y(_2487_));
 sky130_fd_sc_hd__nand2_4 _5911_ (.A(_2485_),
    .B(_2487_),
    .Y(_2488_));
 sky130_fd_sc_hd__nand3b_4 _5912_ (.A_N(_2466_),
    .B(_2482_),
    .C(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__nor2_1 _5913_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .B(_2489_),
    .Y(_2490_));
 sky130_fd_sc_hd__inv_6 _5914_ (.A(_2488_),
    .Y(_2491_));
 sky130_fd_sc_hd__nand2_1 _5915_ (.A(_2491_),
    .B(_2476_),
    .Y(_2492_));
 sky130_fd_sc_hd__inv_2 _5916_ (.A(_2492_),
    .Y(_2493_));
 sky130_fd_sc_hd__nand2_1 _5917_ (.A(_2493_),
    .B(_2466_),
    .Y(_2494_));
 sky130_fd_sc_hd__nor2_1 _5918_ (.A(_2491_),
    .B(_2481_),
    .Y(_2495_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_2495_),
    .B(_2466_),
    .Y(_2496_));
 sky130_fd_sc_hd__o22ai_1 _5920_ (.A1(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .A2(_2494_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .B2(_2496_),
    .Y(_2497_));
 sky130_fd_sc_hd__nor2_1 _5921_ (.A(_2490_),
    .B(_2497_),
    .Y(_2498_));
 sky130_fd_sc_hd__nand3_4 _5922_ (.A(_2464_),
    .B(_2491_),
    .C(_2465_),
    .Y(_2499_));
 sky130_fd_sc_hd__nor2_1 _5923_ (.A(_2477_),
    .B(_2499_),
    .Y(_2500_));
 sky130_fd_sc_hd__nor3_1 _5924_ (.A(_2477_),
    .B(_2491_),
    .C(_2466_),
    .Y(_2501_));
 sky130_fd_sc_hd__inv_2 _5925_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2502_));
 sky130_fd_sc_hd__a22oi_2 _5926_ (.A1(_2500_),
    .A2(_2451_),
    .B1(_2501_),
    .B2(_2502_),
    .Y(_2503_));
 sky130_fd_sc_hd__o21ai_1 _5927_ (.A1(_2481_),
    .A2(_2499_),
    .B1(_2439_),
    .Y(_2504_));
 sky130_fd_sc_hd__nor2_4 _5928_ (.A(_2481_),
    .B(_2499_),
    .Y(_2505_));
 sky130_fd_sc_hd__inv_2 _5929_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2506_));
 sky130_fd_sc_hd__nand2_1 _5930_ (.A(_2505_),
    .B(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__nand2_2 _5931_ (.A(_2504_),
    .B(_2507_),
    .Y(_2508_));
 sky130_fd_sc_hd__nor2_2 _5932_ (.A(_2488_),
    .B(_2481_),
    .Y(_2509_));
 sky130_fd_sc_hd__nand2_1 _5933_ (.A(_2508_),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__nand3_2 _5934_ (.A(_2498_),
    .B(_2503_),
    .C(_2510_),
    .Y(_2511_));
 sky130_fd_sc_hd__buf_6 _5935_ (.A(_2760_),
    .X(_2512_));
 sky130_fd_sc_hd__nand2_2 _5936_ (.A(_2511_),
    .B(_2512_),
    .Y(_2513_));
 sky130_fd_sc_hd__inv_2 _5937_ (.A(_2513_),
    .Y(_2514_));
 sky130_fd_sc_hd__inv_2 _5938_ (.A(_2499_),
    .Y(_2515_));
 sky130_fd_sc_hd__nand2_2 _5939_ (.A(_2515_),
    .B(_2482_),
    .Y(_2516_));
 sky130_fd_sc_hd__nand2_1 _5940_ (.A(_2516_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .Y(_2517_));
 sky130_fd_sc_hd__nand2_1 _5941_ (.A(_2505_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ),
    .Y(_2518_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_2517_),
    .B(_2518_),
    .Y(_2519_));
 sky130_fd_sc_hd__o21ai_1 _5943_ (.A1(_2481_),
    .A2(_2499_),
    .B1(_2441_),
    .Y(_2520_));
 sky130_fd_sc_hd__nand2_1 _5944_ (.A(_2505_),
    .B(_2437_),
    .Y(_2521_));
 sky130_fd_sc_hd__nand2_1 _5945_ (.A(_2520_),
    .B(_2521_),
    .Y(_2522_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(_2519_),
    .B(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__nand2_1 _5947_ (.A(_2516_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2524_));
 sky130_fd_sc_hd__nand2_1 _5948_ (.A(_2505_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ),
    .Y(_2525_));
 sky130_fd_sc_hd__nand2_1 _5949_ (.A(_2524_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_2526_),
    .B(_2508_),
    .Y(_2527_));
 sky130_fd_sc_hd__nand3_1 _5951_ (.A(_2523_),
    .B(_2527_),
    .C(_2509_),
    .Y(_2528_));
 sky130_fd_sc_hd__xnor2_1 _5952_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .Y(_2529_));
 sky130_fd_sc_hd__nand2_1 _5953_ (.A(_2501_),
    .B(_2529_),
    .Y(_2530_));
 sky130_fd_sc_hd__nor2_1 _5954_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2531_));
 sky130_fd_sc_hd__inv_2 _5955_ (.A(_2531_),
    .Y(_2532_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .Y(_2533_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(_2532_),
    .B(_2533_),
    .Y(_2534_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_2500_),
    .B(_2534_),
    .Y(_2535_));
 sky130_fd_sc_hd__nand2_1 _5959_ (.A(_2530_),
    .B(_2535_),
    .Y(_2536_));
 sky130_fd_sc_hd__inv_2 _5960_ (.A(_2489_),
    .Y(_2537_));
 sky130_fd_sc_hd__nand2_1 _5961_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2538_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(_2468_),
    .B(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__nand2_1 _5963_ (.A(_2537_),
    .B(_2539_),
    .Y(_2540_));
 sky130_fd_sc_hd__xor2_1 _5964_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .X(_2541_));
 sky130_fd_sc_hd__nor2_1 _5965_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2542_));
 sky130_fd_sc_hd__inv_2 _5966_ (.A(_2542_),
    .Y(_2543_));
 sky130_fd_sc_hd__nand2_1 _5967_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2544_));
 sky130_fd_sc_hd__nand2_1 _5968_ (.A(_2543_),
    .B(_2544_),
    .Y(_2545_));
 sky130_fd_sc_hd__nand3_1 _5969_ (.A(_2495_),
    .B(_2466_),
    .C(_2545_),
    .Y(_2546_));
 sky130_fd_sc_hd__o21ai_1 _5970_ (.A1(_2541_),
    .A2(_2494_),
    .B1(_2546_),
    .Y(_2547_));
 sky130_fd_sc_hd__inv_2 _5971_ (.A(_2547_),
    .Y(_2548_));
 sky130_fd_sc_hd__nand2_1 _5972_ (.A(_2540_),
    .B(_2548_),
    .Y(_2549_));
 sky130_fd_sc_hd__nor2_1 _5973_ (.A(_2536_),
    .B(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__nand2_1 _5974_ (.A(_2528_),
    .B(_2550_),
    .Y(_2551_));
 sky130_fd_sc_hd__nand2_1 _5975_ (.A(_2551_),
    .B(_2512_),
    .Y(_2552_));
 sky130_fd_sc_hd__nand2_1 _5976_ (.A(_2552_),
    .B(_2513_),
    .Y(_2553_));
 sky130_fd_sc_hd__nor2_2 _5977_ (.A(net17),
    .B(_2759_),
    .Y(_2554_));
 sky130_fd_sc_hd__nand3_1 _5978_ (.A(_2551_),
    .B(_2511_),
    .C(_2512_),
    .Y(_2555_));
 sky130_fd_sc_hd__nand2_1 _5979_ (.A(net17),
    .B(net18),
    .Y(_2556_));
 sky130_fd_sc_hd__inv_2 _5980_ (.A(_2556_),
    .Y(_2557_));
 sky130_fd_sc_hd__and3b_1 _5981_ (.A_N(net21),
    .B(_2557_),
    .C(net20),
    .X(_2558_));
 sky130_fd_sc_hd__inv_2 _5982_ (.A(\egd_top.exp_golomb_decoding.te_range[2] ),
    .Y(_2559_));
 sky130_fd_sc_hd__and2_1 _5983_ (.A(_2558_),
    .B(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__nand2_1 _5984_ (.A(_2466_),
    .B(_2488_),
    .Y(_2561_));
 sky130_fd_sc_hd__o211a_1 _5985_ (.A1(_2479_),
    .A2(_2561_),
    .B1(_2512_),
    .C1(_2480_),
    .X(_2562_));
 sky130_fd_sc_hd__o211a_1 _5986_ (.A1(_2560_),
    .A2(_2511_),
    .B1(_2557_),
    .C1(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__a31o_1 _5987_ (.A1(_2553_),
    .A2(_2554_),
    .A3(_2555_),
    .B1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__a31o_1 _5988_ (.A1(net17),
    .A2(_2759_),
    .A3(_2514_),
    .B1(_2564_),
    .X(net20));
 sky130_fd_sc_hd__a31o_2 _5989_ (.A1(_2558_),
    .A2(net18),
    .A3(_2559_),
    .B1(_2758_),
    .X(_2565_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(_2508_),
    .B(_2522_),
    .Y(_2566_));
 sky130_fd_sc_hd__o21ai_1 _5991_ (.A1(_2481_),
    .A2(_2499_),
    .B1(_2443_),
    .Y(_2567_));
 sky130_fd_sc_hd__nand2_1 _5992_ (.A(_2505_),
    .B(_2439_),
    .Y(_2568_));
 sky130_fd_sc_hd__nand2_1 _5993_ (.A(_2567_),
    .B(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__nand2_1 _5994_ (.A(_2566_),
    .B(_2569_),
    .Y(_2570_));
 sky130_fd_sc_hd__o21ai_1 _5995_ (.A1(_2481_),
    .A2(_2499_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2571_));
 sky130_fd_sc_hd__nand3_1 _5996_ (.A(_2515_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ),
    .C(_2482_),
    .Y(_2572_));
 sky130_fd_sc_hd__nand2_1 _5997_ (.A(_2571_),
    .B(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__nand3_1 _5998_ (.A(_2508_),
    .B(_2522_),
    .C(_2573_),
    .Y(_2574_));
 sky130_fd_sc_hd__nand3_1 _5999_ (.A(_2570_),
    .B(_2574_),
    .C(_2509_),
    .Y(_2575_));
 sky130_fd_sc_hd__nor2_1 _6000_ (.A(_2447_),
    .B(_2467_),
    .Y(_2576_));
 sky130_fd_sc_hd__nor2_1 _6001_ (.A(_2576_),
    .B(_2469_),
    .Y(_2577_));
 sky130_fd_sc_hd__nor2_1 _6002_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ),
    .B(_2532_),
    .Y(_2578_));
 sky130_fd_sc_hd__nor2_1 _6003_ (.A(_2454_),
    .B(_2531_),
    .Y(_2579_));
 sky130_fd_sc_hd__o21ai_1 _6004_ (.A1(_2578_),
    .A2(_2579_),
    .B1(_2500_),
    .Y(_2580_));
 sky130_fd_sc_hd__o21ai_1 _6005_ (.A1(_2577_),
    .A2(_2489_),
    .B1(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__nor2_1 _6006_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ),
    .B(_2542_),
    .Y(_2582_));
 sky130_fd_sc_hd__nor2_1 _6007_ (.A(_2451_),
    .B(_2543_),
    .Y(_2583_));
 sky130_fd_sc_hd__and2_1 _6008_ (.A(_2455_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ),
    .X(_2584_));
 sky130_fd_sc_hd__o21bai_1 _6009_ (.A1(_2456_),
    .A2(_2584_),
    .B1_N(_2494_),
    .Y(_2585_));
 sky130_fd_sc_hd__o31ai_1 _6010_ (.A1(_2582_),
    .A2(_2583_),
    .A3(_2496_),
    .B1(_2585_),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_1 _6011_ (.A(_2581_),
    .B(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__nand2_1 _6012_ (.A(_2575_),
    .B(_2587_),
    .Y(_2588_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(_2588_),
    .B(_2512_),
    .Y(_2589_));
 sky130_fd_sc_hd__nand2_1 _6014_ (.A(_2589_),
    .B(_2552_),
    .Y(_2590_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(_2590_),
    .B(_2554_),
    .Y(_2591_));
 sky130_fd_sc_hd__a31o_1 _6016_ (.A1(_2562_),
    .A2(_2551_),
    .A3(_2588_),
    .B1(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__o21ai_2 _6017_ (.A1(_2552_),
    .A2(_2565_),
    .B1(_2592_),
    .Y(net21));
 sky130_fd_sc_hd__o21ai_1 _6018_ (.A1(_2552_),
    .A2(_2589_),
    .B1(_2514_),
    .Y(_2593_));
 sky130_fd_sc_hd__nand2_1 _6019_ (.A(_2593_),
    .B(_2590_),
    .Y(_2594_));
 sky130_fd_sc_hd__nor2_1 _6020_ (.A(_2519_),
    .B(_2526_),
    .Y(_2595_));
 sky130_fd_sc_hd__nand2_1 _6021_ (.A(_2516_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2596_));
 sky130_fd_sc_hd__nand2_1 _6022_ (.A(_2505_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ),
    .Y(_2597_));
 sky130_fd_sc_hd__nand2_1 _6023_ (.A(_2596_),
    .B(_2597_),
    .Y(_2598_));
 sky130_fd_sc_hd__nand3_1 _6024_ (.A(_2595_),
    .B(_2569_),
    .C(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__nand3_1 _6025_ (.A(_2508_),
    .B(_2522_),
    .C(_2569_),
    .Y(_2600_));
 sky130_fd_sc_hd__nand2_1 _6026_ (.A(_2516_),
    .B(_2445_),
    .Y(_2601_));
 sky130_fd_sc_hd__nand2_1 _6027_ (.A(_2505_),
    .B(_2441_),
    .Y(_2602_));
 sky130_fd_sc_hd__nand2_1 _6028_ (.A(_2601_),
    .B(_2602_),
    .Y(_2603_));
 sky130_fd_sc_hd__nand2_1 _6029_ (.A(_2600_),
    .B(_2603_),
    .Y(_2604_));
 sky130_fd_sc_hd__nand3_1 _6030_ (.A(_2599_),
    .B(_2509_),
    .C(_2604_),
    .Y(_2605_));
 sky130_fd_sc_hd__nand2_1 _6031_ (.A(_2543_),
    .B(_2457_),
    .Y(_2606_));
 sky130_fd_sc_hd__o21ai_1 _6032_ (.A1(_2543_),
    .A2(_2534_),
    .B1(_2606_),
    .Y(_2607_));
 sky130_fd_sc_hd__nor2_1 _6033_ (.A(_2468_),
    .B(_2543_),
    .Y(_2608_));
 sky130_fd_sc_hd__nor2_1 _6034_ (.A(_2449_),
    .B(_2469_),
    .Y(_2609_));
 sky130_fd_sc_hd__nor2_1 _6035_ (.A(_2608_),
    .B(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__nor2_1 _6036_ (.A(_2455_),
    .B(_2532_),
    .Y(_2611_));
 sky130_fd_sc_hd__nor2_1 _6037_ (.A(_2453_),
    .B(_2578_),
    .Y(_2612_));
 sky130_fd_sc_hd__o21ai_1 _6038_ (.A1(_2611_),
    .A2(_2612_),
    .B1(_2500_),
    .Y(_2613_));
 sky130_fd_sc_hd__o221a_1 _6039_ (.A1(_2496_),
    .A2(_2607_),
    .B1(_2610_),
    .B2(_2489_),
    .C1(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__inv_2 _6040_ (.A(_2760_),
    .Y(_2615_));
 sky130_fd_sc_hd__a21oi_1 _6041_ (.A1(_2605_),
    .A2(_2614_),
    .B1(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_2594_),
    .B(_2616_),
    .Y(_2617_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(_2605_),
    .B(_2614_),
    .Y(_2618_));
 sky130_fd_sc_hd__nand2_1 _6044_ (.A(_2618_),
    .B(_2512_),
    .Y(_2619_));
 sky130_fd_sc_hd__nand3_1 _6045_ (.A(_2593_),
    .B(_2590_),
    .C(_2619_),
    .Y(_2620_));
 sky130_fd_sc_hd__nand2_1 _6046_ (.A(_2617_),
    .B(_2620_),
    .Y(_2621_));
 sky130_fd_sc_hd__nand2_1 _6047_ (.A(_2621_),
    .B(_2554_),
    .Y(_2622_));
 sky130_fd_sc_hd__or2_1 _6048_ (.A(_2565_),
    .B(_2589_),
    .X(_2623_));
 sky130_fd_sc_hd__nand2_1 _6049_ (.A(net20),
    .B(net21),
    .Y(_2624_));
 sky130_fd_sc_hd__a21oi_1 _6050_ (.A1(_2622_),
    .A2(_2623_),
    .B1(_2624_),
    .Y(_2625_));
 sky130_fd_sc_hd__nand3_1 _6051_ (.A(_2622_),
    .B(_2624_),
    .C(_2623_),
    .Y(_2626_));
 sky130_fd_sc_hd__nand2_1 _6052_ (.A(_2626_),
    .B(_2557_),
    .Y(_2627_));
 sky130_fd_sc_hd__nor2_1 _6053_ (.A(_2625_),
    .B(_2627_),
    .Y(\egd_top.exp_golomb_decoding.te_range[2] ));
 sky130_fd_sc_hd__or3_1 _6054_ (.A(_2615_),
    .B(_2560_),
    .C(_2478_),
    .X(_2628_));
 sky130_fd_sc_hd__inv_2 _6055_ (.A(_2628_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[3] ));
 sky130_fd_sc_hd__or3_1 _6056_ (.A(_2615_),
    .B(_2560_),
    .C(_2488_),
    .X(_2629_));
 sky130_fd_sc_hd__inv_2 _6057_ (.A(_2629_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[2] ));
 sky130_fd_sc_hd__or3_1 _6058_ (.A(_2615_),
    .B(_2560_),
    .C(_2466_),
    .X(_2630_));
 sky130_fd_sc_hd__inv_2 _6059_ (.A(_2630_),
    .Y(\egd_top.BitStream_buffer.exp_golomb_len[1] ));
 sky130_fd_sc_hd__nand2_1 _6060_ (.A(_2622_),
    .B(_2623_),
    .Y(net22));
 sky130_fd_sc_hd__nand2_1 _6061_ (.A(_2603_),
    .B(_2569_),
    .Y(_2631_));
 sky130_fd_sc_hd__o21ai_1 _6062_ (.A1(_2481_),
    .A2(_2499_),
    .B1(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ),
    .Y(_2632_));
 sky130_fd_sc_hd__nand2_1 _6063_ (.A(_2505_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ),
    .Y(_2633_));
 sky130_fd_sc_hd__nand2_1 _6064_ (.A(_2632_),
    .B(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__inv_2 _6065_ (.A(_2634_),
    .Y(_2635_));
 sky130_fd_sc_hd__o21ai_1 _6066_ (.A1(_2566_),
    .A2(_2631_),
    .B1(_2635_),
    .Y(_2636_));
 sky130_fd_sc_hd__nor2_1 _6067_ (.A(_2566_),
    .B(_2631_),
    .Y(_2637_));
 sky130_fd_sc_hd__nand2_1 _6068_ (.A(_2637_),
    .B(_2634_),
    .Y(_2638_));
 sky130_fd_sc_hd__nand3_1 _6069_ (.A(_2636_),
    .B(_2638_),
    .C(_2509_),
    .Y(_2639_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_2542_),
    .B(_2531_),
    .Y(_2640_));
 sky130_fd_sc_hd__and2_1 _6071_ (.A(_2640_),
    .B(_2454_),
    .X(_2641_));
 sky130_fd_sc_hd__nor2_1 _6072_ (.A(_2454_),
    .B(_2640_),
    .Y(_2642_));
 sky130_fd_sc_hd__xor2_1 _6073_ (.A(_2451_),
    .B(_2608_),
    .X(_2643_));
 sky130_fd_sc_hd__o32a_1 _6074_ (.A1(_2641_),
    .A2(_2642_),
    .A3(_2496_),
    .B1(_2489_),
    .B2(_2643_),
    .X(_2644_));
 sky130_fd_sc_hd__nand2_1 _6075_ (.A(_2639_),
    .B(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__nand2_1 _6076_ (.A(_2645_),
    .B(_2512_),
    .Y(_2646_));
 sky130_fd_sc_hd__nor2_1 _6077_ (.A(_2555_),
    .B(_2589_),
    .Y(_2647_));
 sky130_fd_sc_hd__nand2_2 _6078_ (.A(_2616_),
    .B(_2647_),
    .Y(_2648_));
 sky130_fd_sc_hd__nor2_1 _6079_ (.A(_2646_),
    .B(_2648_),
    .Y(_2649_));
 sky130_fd_sc_hd__a21oi_2 _6080_ (.A1(_2639_),
    .A2(_2644_),
    .B1(_2615_),
    .Y(_2650_));
 sky130_fd_sc_hd__inv_2 _6081_ (.A(_2648_),
    .Y(_2651_));
 sky130_fd_sc_hd__nor2_1 _6082_ (.A(_2650_),
    .B(_2651_),
    .Y(_2652_));
 sky130_fd_sc_hd__o21ai_1 _6083_ (.A1(_2649_),
    .A2(_2652_),
    .B1(_2514_),
    .Y(_2653_));
 sky130_fd_sc_hd__o21bai_1 _6084_ (.A1(_2551_),
    .A2(_2588_),
    .B1_N(_2615_),
    .Y(_2654_));
 sky130_fd_sc_hd__nand2_1 _6085_ (.A(_2654_),
    .B(_2619_),
    .Y(_2655_));
 sky130_fd_sc_hd__nor2_2 _6086_ (.A(_2650_),
    .B(_2655_),
    .Y(_2656_));
 sky130_fd_sc_hd__and2_1 _6087_ (.A(_2655_),
    .B(_2650_),
    .X(_2657_));
 sky130_fd_sc_hd__o21ai_1 _6088_ (.A1(_2656_),
    .A2(_2657_),
    .B1(_2513_),
    .Y(_2658_));
 sky130_fd_sc_hd__nand3_1 _6089_ (.A(_2653_),
    .B(_2554_),
    .C(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__o21ai_2 _6090_ (.A1(_2619_),
    .A2(_2565_),
    .B1(_2659_),
    .Y(net23));
 sky130_fd_sc_hd__o21ai_1 _6091_ (.A1(_2646_),
    .A2(_2648_),
    .B1(_2514_),
    .Y(_2660_));
 sky130_fd_sc_hd__nand2_1 _6092_ (.A(_2656_),
    .B(_2513_),
    .Y(_2661_));
 sky130_fd_sc_hd__nand2_1 _6093_ (.A(_2660_),
    .B(_2661_),
    .Y(_2662_));
 sky130_fd_sc_hd__nor2_1 _6094_ (.A(_2573_),
    .B(_2598_),
    .Y(_2663_));
 sky130_fd_sc_hd__nand3_1 _6095_ (.A(_2595_),
    .B(_2663_),
    .C(_2635_),
    .Y(_2664_));
 sky130_fd_sc_hd__nand2_1 _6096_ (.A(_2516_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ),
    .Y(_2665_));
 sky130_fd_sc_hd__nand2_1 _6097_ (.A(_2505_),
    .B(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ),
    .Y(_2666_));
 sky130_fd_sc_hd__nand2_1 _6098_ (.A(_2665_),
    .B(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__inv_2 _6099_ (.A(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__nand2_1 _6100_ (.A(_2664_),
    .B(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__nand3_1 _6101_ (.A(_2637_),
    .B(_2635_),
    .C(_2667_),
    .Y(_2670_));
 sky130_fd_sc_hd__nand3_1 _6102_ (.A(_2669_),
    .B(_2670_),
    .C(_2509_),
    .Y(_2671_));
 sky130_fd_sc_hd__nor2_1 _6103_ (.A(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ),
    .B(_2608_),
    .Y(_2672_));
 sky130_fd_sc_hd__a311o_1 _6104_ (.A1(_2532_),
    .A2(_2608_),
    .A3(_2533_),
    .B1(_2672_),
    .C1(_2489_),
    .X(_2673_));
 sky130_fd_sc_hd__nand2_1 _6105_ (.A(_2671_),
    .B(_2673_),
    .Y(_2674_));
 sky130_fd_sc_hd__nand2_1 _6106_ (.A(_2674_),
    .B(_2512_),
    .Y(_2675_));
 sky130_fd_sc_hd__nand2_1 _6107_ (.A(_2662_),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__inv_2 _6108_ (.A(_2675_),
    .Y(_2677_));
 sky130_fd_sc_hd__nand3_1 _6109_ (.A(_2660_),
    .B(_2677_),
    .C(_2661_),
    .Y(_2678_));
 sky130_fd_sc_hd__nand3_1 _6110_ (.A(_2676_),
    .B(_2554_),
    .C(_2678_),
    .Y(_2679_));
 sky130_fd_sc_hd__o21ai_2 _6111_ (.A1(_2646_),
    .A2(_2565_),
    .B1(_2679_),
    .Y(net24));
 sky130_fd_sc_hd__nand2_1 _6112_ (.A(_2656_),
    .B(_2675_),
    .Y(_2680_));
 sky130_fd_sc_hd__inv_2 _6113_ (.A(_2509_),
    .Y(_2681_));
 sky130_fd_sc_hd__nor2_1 _6114_ (.A(_2634_),
    .B(_2667_),
    .Y(_2682_));
 sky130_fd_sc_hd__nand3_1 _6115_ (.A(_2595_),
    .B(_2663_),
    .C(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__o21ai_2 _6116_ (.A1(_2447_),
    .A2(_2516_),
    .B1(_2451_),
    .Y(_2684_));
 sky130_fd_sc_hd__inv_2 _6117_ (.A(_2684_),
    .Y(_2685_));
 sky130_fd_sc_hd__nand2_1 _6118_ (.A(_2683_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__nand3_1 _6119_ (.A(_2637_),
    .B(_2682_),
    .C(_2684_),
    .Y(_2687_));
 sky130_fd_sc_hd__nand2_1 _6120_ (.A(_2686_),
    .B(_2687_),
    .Y(_2688_));
 sky130_fd_sc_hd__nor2_1 _6121_ (.A(_2681_),
    .B(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__nand2_1 _6122_ (.A(_2689_),
    .B(_2512_),
    .Y(_2690_));
 sky130_fd_sc_hd__inv_2 _6123_ (.A(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__nand2_1 _6124_ (.A(_2680_),
    .B(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__o21ai_1 _6125_ (.A1(_2689_),
    .A2(_2674_),
    .B1(_2512_),
    .Y(_2693_));
 sky130_fd_sc_hd__nand2_1 _6126_ (.A(_2693_),
    .B(_2656_),
    .Y(_2694_));
 sky130_fd_sc_hd__nand3_1 _6127_ (.A(_2692_),
    .B(_2513_),
    .C(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__nand3_1 _6128_ (.A(_2649_),
    .B(_2691_),
    .C(_2677_),
    .Y(_2696_));
 sky130_fd_sc_hd__nand3_1 _6129_ (.A(_2674_),
    .B(_2512_),
    .C(_2645_),
    .Y(_2697_));
 sky130_fd_sc_hd__o21ai_1 _6130_ (.A1(_2648_),
    .A2(_2697_),
    .B1(_2690_),
    .Y(_2698_));
 sky130_fd_sc_hd__nand3_1 _6131_ (.A(_2696_),
    .B(_2698_),
    .C(_2514_),
    .Y(_2699_));
 sky130_fd_sc_hd__nand2_1 _6132_ (.A(_2695_),
    .B(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__nand2_1 _6133_ (.A(_2700_),
    .B(_2554_),
    .Y(_2701_));
 sky130_fd_sc_hd__inv_2 _6134_ (.A(_2565_),
    .Y(_2702_));
 sky130_fd_sc_hd__nand2_1 _6135_ (.A(_2677_),
    .B(_2702_),
    .Y(_2703_));
 sky130_fd_sc_hd__nand2_1 _6136_ (.A(_2701_),
    .B(_2703_),
    .Y(net25));
 sky130_fd_sc_hd__or2_1 _6137_ (.A(_2684_),
    .B(_2683_),
    .X(_2704_));
 sky130_fd_sc_hd__nand3_1 _6138_ (.A(_2704_),
    .B(_2512_),
    .C(_2505_),
    .Y(_2705_));
 sky130_fd_sc_hd__inv_2 _6139_ (.A(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__nand2_1 _6140_ (.A(_2694_),
    .B(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__nand3_1 _6141_ (.A(_2704_),
    .B(_2505_),
    .C(_2562_),
    .Y(_2708_));
 sky130_fd_sc_hd__nand3_1 _6142_ (.A(_2693_),
    .B(_2656_),
    .C(_2708_),
    .Y(_2709_));
 sky130_fd_sc_hd__nand2_1 _6143_ (.A(_2707_),
    .B(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__nand2_1 _6144_ (.A(_2710_),
    .B(_2513_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand3b_1 _6145_ (.A_N(_2697_),
    .B(_2691_),
    .C(_2651_),
    .Y(_2712_));
 sky130_fd_sc_hd__nand3_1 _6146_ (.A(_2712_),
    .B(_2514_),
    .C(_2705_),
    .Y(_2713_));
 sky130_fd_sc_hd__nand3_1 _6147_ (.A(_2711_),
    .B(_2554_),
    .C(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__nand2_1 _6148_ (.A(_2691_),
    .B(_2702_),
    .Y(_2715_));
 sky130_fd_sc_hd__nand2_1 _6149_ (.A(_2714_),
    .B(_2715_),
    .Y(net26));
 sky130_fd_sc_hd__nor2_1 _6150_ (.A(_2565_),
    .B(_2708_),
    .Y(_2716_));
 sky130_fd_sc_hd__a31o_1 _6151_ (.A1(_2562_),
    .A2(_2513_),
    .A3(_2554_),
    .B1(_2716_),
    .X(net27));
 sky130_fd_sc_hd__buf_1 _6152_ (.A(clknet_1_0__leaf_wb_clk_i),
    .X(_2717_));
 sky130_fd_sc_hd__buf_1 _6153_ (.A(clknet_1_1__leaf__2717_),
    .X(_2718_));
 sky130_fd_sc_hd__inv_2 _6154__25 (.A(clknet_1_0__leaf__2718_),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _6155__26 (.A(clknet_1_0__leaf__2718_),
    .Y(net78));
 sky130_fd_sc_hd__inv_2 _6156__27 (.A(clknet_1_0__leaf__2718_),
    .Y(net79));
 sky130_fd_sc_hd__inv_2 _6157__28 (.A(clknet_1_0__leaf__2718_),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _6158__29 (.A(clknet_1_0__leaf__2718_),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _6159__30 (.A(clknet_1_1__leaf__2718_),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _6160__31 (.A(clknet_1_1__leaf__2718_),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _6161__32 (.A(clknet_1_1__leaf__2718_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _6162__33 (.A(clknet_1_1__leaf__2718_),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _6163__34 (.A(clknet_1_1__leaf__2718_),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _6164__35 (.A(clknet_1_1__leaf__2718_),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _6165__36 (.A(clknet_1_1__leaf__2718_),
    .Y(net88));
 sky130_fd_sc_hd__buf_1 _6166_ (.A(clknet_1_0__leaf__2717_),
    .X(_2719_));
 sky130_fd_sc_hd__inv_2 _6167__37 (.A(clknet_1_1__leaf__2719_),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _6168__38 (.A(clknet_1_1__leaf__2719_),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _6169__39 (.A(clknet_1_1__leaf__2719_),
    .Y(net91));
 sky130_fd_sc_hd__inv_2 _6170__40 (.A(clknet_1_1__leaf__2719_),
    .Y(net92));
 sky130_fd_sc_hd__inv_2 _6171__41 (.A(clknet_1_0__leaf__2719_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _6172__42 (.A(clknet_1_0__leaf__2719_),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _6173__43 (.A(clknet_1_0__leaf__2719_),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _6174__44 (.A(clknet_1_0__leaf__2719_),
    .Y(net96));
 sky130_fd_sc_hd__inv_2 _6175__45 (.A(clknet_1_0__leaf__2719_),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _6176__46 (.A(clknet_1_0__leaf__2719_),
    .Y(net98));
 sky130_fd_sc_hd__inv_2 _6177__47 (.A(clknet_1_0__leaf__2719_),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _6178__48 (.A(clknet_1_1__leaf__2719_),
    .Y(net100));
 sky130_fd_sc_hd__buf_1 _6179_ (.A(clknet_1_0__leaf__2717_),
    .X(_2720_));
 sky130_fd_sc_hd__inv_2 _6180__49 (.A(clknet_1_1__leaf__2720_),
    .Y(net101));
 sky130_fd_sc_hd__inv_2 _6181__50 (.A(clknet_1_1__leaf__2720_),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _6182__51 (.A(clknet_1_1__leaf__2720_),
    .Y(net103));
 sky130_fd_sc_hd__inv_2 _6183__52 (.A(clknet_1_1__leaf__2720_),
    .Y(net104));
 sky130_fd_sc_hd__inv_2 _6184__53 (.A(clknet_1_1__leaf__2720_),
    .Y(net105));
 sky130_fd_sc_hd__inv_2 _6185__54 (.A(clknet_1_0__leaf__2720_),
    .Y(net106));
 sky130_fd_sc_hd__inv_2 _6186__55 (.A(clknet_1_1__leaf__2720_),
    .Y(net107));
 sky130_fd_sc_hd__inv_2 _6187__56 (.A(clknet_1_0__leaf__2720_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _6188__57 (.A(clknet_1_0__leaf__2720_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _6189__58 (.A(clknet_1_0__leaf__2720_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _6190__59 (.A(clknet_1_0__leaf__2720_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _6191__60 (.A(clknet_1_0__leaf__2720_),
    .Y(net112));
 sky130_fd_sc_hd__buf_1 _6192_ (.A(clknet_1_0__leaf__2717_),
    .X(_2721_));
 sky130_fd_sc_hd__inv_2 _6193__61 (.A(clknet_1_0__leaf__2721_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _6194__62 (.A(clknet_1_0__leaf__2721_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _6195__63 (.A(clknet_1_0__leaf__2721_),
    .Y(net115));
 sky130_fd_sc_hd__inv_2 _6196__64 (.A(clknet_1_0__leaf__2721_),
    .Y(net116));
 sky130_fd_sc_hd__inv_2 _6197__65 (.A(clknet_1_0__leaf__2721_),
    .Y(net117));
 sky130_fd_sc_hd__inv_2 _6198__66 (.A(clknet_1_0__leaf__2721_),
    .Y(net118));
 sky130_fd_sc_hd__inv_2 _6199__67 (.A(clknet_1_1__leaf__2721_),
    .Y(net119));
 sky130_fd_sc_hd__inv_2 _6200__68 (.A(clknet_1_1__leaf__2721_),
    .Y(net120));
 sky130_fd_sc_hd__inv_2 _6201__69 (.A(clknet_1_1__leaf__2721_),
    .Y(net121));
 sky130_fd_sc_hd__inv_2 _6202__70 (.A(clknet_1_1__leaf__2721_),
    .Y(net122));
 sky130_fd_sc_hd__inv_2 _6203__71 (.A(clknet_1_1__leaf__2721_),
    .Y(net123));
 sky130_fd_sc_hd__inv_2 _6204__72 (.A(clknet_1_1__leaf__2721_),
    .Y(net124));
 sky130_fd_sc_hd__buf_1 _6205_ (.A(clknet_1_1__leaf__2717_),
    .X(_2722_));
 sky130_fd_sc_hd__inv_2 _6206__73 (.A(clknet_1_0__leaf__2722_),
    .Y(net125));
 sky130_fd_sc_hd__inv_2 _6207__74 (.A(clknet_1_0__leaf__2722_),
    .Y(net126));
 sky130_fd_sc_hd__inv_2 _6208__75 (.A(clknet_1_0__leaf__2722_),
    .Y(net127));
 sky130_fd_sc_hd__inv_2 _6209__76 (.A(clknet_1_1__leaf__2722_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _6210__77 (.A(clknet_1_1__leaf__2722_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _6211__78 (.A(clknet_1_1__leaf__2722_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _6212__79 (.A(clknet_1_1__leaf__2722_),
    .Y(net131));
 sky130_fd_sc_hd__inv_2 _6213__80 (.A(clknet_1_1__leaf__2722_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _6214__81 (.A(clknet_1_1__leaf__2722_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _6215__82 (.A(clknet_1_0__leaf__2722_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _6216__83 (.A(clknet_1_0__leaf__2722_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _6217__84 (.A(clknet_1_0__leaf__2722_),
    .Y(net136));
 sky130_fd_sc_hd__buf_1 _6218_ (.A(clknet_1_1__leaf__2717_),
    .X(_2723_));
 sky130_fd_sc_hd__inv_2 _6219__85 (.A(clknet_1_0__leaf__2723_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _6220__86 (.A(clknet_1_0__leaf__2723_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _6221__87 (.A(clknet_1_0__leaf__2723_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _6222__88 (.A(clknet_1_0__leaf__2723_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _6223__89 (.A(clknet_1_0__leaf__2723_),
    .Y(net141));
 sky130_fd_sc_hd__inv_2 _6224__90 (.A(clknet_1_1__leaf__2723_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _6225__91 (.A(clknet_1_1__leaf__2723_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _6226__92 (.A(clknet_1_1__leaf__2723_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _6227__93 (.A(clknet_1_1__leaf__2723_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _6228__94 (.A(clknet_1_1__leaf__2723_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _6229__95 (.A(clknet_1_1__leaf__2723_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _6230__96 (.A(clknet_1_1__leaf__2723_),
    .Y(net148));
 sky130_fd_sc_hd__buf_1 _6231_ (.A(clknet_1_1__leaf__2717_),
    .X(_2724_));
 sky130_fd_sc_hd__inv_2 _6232__97 (.A(clknet_1_1__leaf__2724_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _6233__98 (.A(clknet_1_1__leaf__2724_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _6234__99 (.A(clknet_1_0__leaf__2724_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _6235__100 (.A(clknet_1_0__leaf__2724_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _6236__101 (.A(clknet_1_0__leaf__2724_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _6237__102 (.A(clknet_1_0__leaf__2724_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _6238__103 (.A(clknet_1_0__leaf__2724_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _6239__104 (.A(clknet_1_0__leaf__2724_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _6240__105 (.A(clknet_1_1__leaf__2724_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _6241__106 (.A(clknet_1_1__leaf__2724_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _6242__107 (.A(clknet_1_1__leaf__2724_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _6243__108 (.A(clknet_1_1__leaf__2724_),
    .Y(net160));
 sky130_fd_sc_hd__buf_1 _6244_ (.A(clknet_1_1__leaf__2717_),
    .X(_2725_));
 sky130_fd_sc_hd__inv_2 _6245__109 (.A(clknet_1_1__leaf__2725_),
    .Y(net161));
 sky130_fd_sc_hd__inv_2 _6246__110 (.A(clknet_1_1__leaf__2725_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _6247__111 (.A(clknet_1_1__leaf__2725_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _6248__112 (.A(clknet_1_1__leaf__2725_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _6249__113 (.A(clknet_1_1__leaf__2725_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _6250__114 (.A(clknet_1_1__leaf__2725_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _6251__115 (.A(clknet_1_0__leaf__2725_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _6252__116 (.A(clknet_1_0__leaf__2725_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _6253__117 (.A(clknet_1_0__leaf__2725_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _6254__118 (.A(clknet_1_0__leaf__2725_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _6255__119 (.A(clknet_1_0__leaf__2725_),
    .Y(net171));
 sky130_fd_sc_hd__inv_2 _6256__120 (.A(clknet_1_1__leaf__2725_),
    .Y(net172));
 sky130_fd_sc_hd__buf_1 _6257_ (.A(clknet_1_0__leaf__2717_),
    .X(_2726_));
 sky130_fd_sc_hd__inv_2 _6258__121 (.A(clknet_1_0__leaf__2726_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _6259__122 (.A(clknet_1_1__leaf__2726_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _6260__123 (.A(clknet_1_1__leaf__2726_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _6261__124 (.A(clknet_1_1__leaf__2726_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _6262__125 (.A(clknet_1_1__leaf__2726_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _6263__126 (.A(clknet_1_1__leaf__2726_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _6264__127 (.A(clknet_1_1__leaf__2726_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _6265__128 (.A(clknet_1_1__leaf__2726_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _6266__129 (.A(clknet_1_0__leaf__2726_),
    .Y(net181));
 sky130_fd_sc_hd__inv_2 _6267__130 (.A(clknet_1_0__leaf__2726_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _6268__131 (.A(clknet_1_0__leaf__2726_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _6269__132 (.A(clknet_1_0__leaf__2726_),
    .Y(net184));
 sky130_fd_sc_hd__buf_1 _6270_ (.A(clknet_1_0__leaf__2717_),
    .X(_2727_));
 sky130_fd_sc_hd__inv_2 _6271__133 (.A(clknet_1_0__leaf__2727_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _6272__134 (.A(clknet_1_1__leaf__2727_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _6273__135 (.A(clknet_1_1__leaf__2727_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _6274__136 (.A(clknet_1_0__leaf__2727_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _6275__137 (.A(clknet_1_0__leaf__2727_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _6276__138 (.A(clknet_1_0__leaf__2727_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _6277__139 (.A(clknet_1_1__leaf__2727_),
    .Y(net191));
 sky130_fd_sc_hd__inv_2 _6278__140 (.A(clknet_1_0__leaf__2727_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _6279__141 (.A(clknet_1_0__leaf__2727_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _6280__142 (.A(clknet_1_0__leaf__2727_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _6281__143 (.A(clknet_1_1__leaf__2727_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _6282__144 (.A(clknet_1_1__leaf__2727_),
    .Y(net196));
 sky130_fd_sc_hd__buf_1 _6283_ (.A(clknet_1_0__leaf__2717_),
    .X(_2728_));
 sky130_fd_sc_hd__inv_2 _6284__145 (.A(clknet_1_1__leaf__2728_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _6285__146 (.A(clknet_1_1__leaf__2728_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _6286__147 (.A(clknet_1_0__leaf__2728_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _6287__148 (.A(clknet_1_0__leaf__2728_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _6288__149 (.A(clknet_1_0__leaf__2728_),
    .Y(net201));
 sky130_fd_sc_hd__inv_2 _6289__150 (.A(clknet_1_0__leaf__2728_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _6290__151 (.A(clknet_1_0__leaf__2728_),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _6291__152 (.A(clknet_1_0__leaf__2728_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _6292__153 (.A(clknet_1_1__leaf__2728_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _6293__154 (.A(clknet_1_1__leaf__2728_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _6294__155 (.A(clknet_1_1__leaf__2728_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _6295__156 (.A(clknet_1_1__leaf__2728_),
    .Y(net208));
 sky130_fd_sc_hd__buf_1 _6296_ (.A(clknet_1_0__leaf__2717_),
    .X(_2729_));
 sky130_fd_sc_hd__inv_2 _6297__157 (.A(clknet_1_0__leaf__2729_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _6298__158 (.A(clknet_1_0__leaf__2729_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _6299__159 (.A(clknet_1_0__leaf__2729_),
    .Y(net211));
 sky130_fd_sc_hd__inv_2 _6300__160 (.A(clknet_1_0__leaf__2729_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _6301__161 (.A(clknet_1_0__leaf__2729_),
    .Y(net213));
 sky130_fd_sc_hd__inv_2 _6302__162 (.A(clknet_1_0__leaf__2729_),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _6303__163 (.A(clknet_1_1__leaf__2729_),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _6304__164 (.A(clknet_1_1__leaf__2729_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _6305__165 (.A(clknet_1_1__leaf__2729_),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _6306__166 (.A(clknet_1_1__leaf__2729_),
    .Y(net218));
 sky130_fd_sc_hd__inv_2 _6307__167 (.A(clknet_1_1__leaf__2729_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _6308__168 (.A(clknet_1_1__leaf__2729_),
    .Y(net220));
 sky130_fd_sc_hd__buf_1 _6309_ (.A(clknet_1_1__leaf_wb_clk_i),
    .X(_2730_));
 sky130_fd_sc_hd__inv_2 _6310__1 (.A(clknet_1_1__leaf__2730_),
    .Y(net53));
 sky130_fd_sc_hd__inv_2 _6311__2 (.A(clknet_1_1__leaf__2730_),
    .Y(net54));
 sky130_fd_sc_hd__inv_2 _6312__3 (.A(clknet_1_1__leaf__2730_),
    .Y(net55));
 sky130_fd_sc_hd__inv_2 _6313__4 (.A(clknet_1_1__leaf__2730_),
    .Y(net56));
 sky130_fd_sc_hd__inv_2 _6314__5 (.A(clknet_1_1__leaf__2730_),
    .Y(net57));
 sky130_fd_sc_hd__inv_2 _6315__6 (.A(clknet_1_1__leaf__2730_),
    .Y(net58));
 sky130_fd_sc_hd__inv_2 _6316__7 (.A(clknet_1_1__leaf__2730_),
    .Y(net59));
 sky130_fd_sc_hd__inv_2 _6317__8 (.A(clknet_1_0__leaf__2730_),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 _6318__9 (.A(clknet_1_0__leaf__2730_),
    .Y(net61));
 sky130_fd_sc_hd__inv_2 _6319__10 (.A(clknet_1_0__leaf__2730_),
    .Y(net62));
 sky130_fd_sc_hd__inv_2 _6320__11 (.A(clknet_1_0__leaf__2730_),
    .Y(net63));
 sky130_fd_sc_hd__inv_2 _6321__12 (.A(clknet_1_0__leaf__2730_),
    .Y(net64));
 sky130_fd_sc_hd__buf_1 _6322_ (.A(clknet_1_0__leaf_wb_clk_i),
    .X(_2731_));
 sky130_fd_sc_hd__inv_2 _6323__13 (.A(clknet_1_0__leaf__2731_),
    .Y(net65));
 sky130_fd_sc_hd__inv_2 _6324__14 (.A(clknet_1_1__leaf__2731_),
    .Y(net66));
 sky130_fd_sc_hd__inv_2 _6325__15 (.A(clknet_1_1__leaf__2731_),
    .Y(net67));
 sky130_fd_sc_hd__inv_2 _6326__16 (.A(clknet_1_1__leaf__2731_),
    .Y(net68));
 sky130_fd_sc_hd__inv_2 _6327__17 (.A(clknet_1_1__leaf__2731_),
    .Y(net69));
 sky130_fd_sc_hd__inv_2 _6328__18 (.A(clknet_1_1__leaf__2731_),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _6329__19 (.A(clknet_1_1__leaf__2731_),
    .Y(net71));
 sky130_fd_sc_hd__inv_2 _6330__20 (.A(clknet_1_0__leaf__2731_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _6331__21 (.A(clknet_1_0__leaf__2731_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _6332__22 (.A(clknet_1_0__leaf__2731_),
    .Y(net74));
 sky130_fd_sc_hd__inv_2 _6333__23 (.A(clknet_1_0__leaf__2731_),
    .Y(net75));
 sky130_fd_sc_hd__inv_2 _6334__24 (.A(clknet_1_0__leaf__2731_),
    .Y(net76));
 sky130_fd_sc_hd__dfrtp_1 _6335_ (.CLK(net77),
    .D(_0168_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[95] ));
 sky130_fd_sc_hd__dfrtp_4 _6336_ (.CLK(net78),
    .D(_0169_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[94] ));
 sky130_fd_sc_hd__dfrtp_2 _6337_ (.CLK(net79),
    .D(_0170_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[93] ));
 sky130_fd_sc_hd__dfrtp_2 _6338_ (.CLK(net80),
    .D(_0171_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[92] ));
 sky130_fd_sc_hd__dfrtp_4 _6339_ (.CLK(net81),
    .D(_0172_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[91] ));
 sky130_fd_sc_hd__dfrtp_4 _6340_ (.CLK(net82),
    .D(_0173_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[90] ));
 sky130_fd_sc_hd__dfrtp_4 _6341_ (.CLK(net83),
    .D(_0174_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[89] ));
 sky130_fd_sc_hd__dfrtp_4 _6342_ (.CLK(net84),
    .D(_0175_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[88] ));
 sky130_fd_sc_hd__dfrtp_2 _6343_ (.CLK(net85),
    .D(_0176_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[87] ));
 sky130_fd_sc_hd__dfrtp_4 _6344_ (.CLK(net86),
    .D(_0177_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[86] ));
 sky130_fd_sc_hd__dfrtp_4 _6345_ (.CLK(net87),
    .D(_0178_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[85] ));
 sky130_fd_sc_hd__dfrtp_4 _6346_ (.CLK(net88),
    .D(_0179_),
    .RESET_B(net51),
    .Q(\egd_top.BitStream_buffer.BS_buffer[84] ));
 sky130_fd_sc_hd__dfrtp_4 _6347_ (.CLK(net89),
    .D(_0180_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[83] ));
 sky130_fd_sc_hd__dfrtp_4 _6348_ (.CLK(net90),
    .D(_0181_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[82] ));
 sky130_fd_sc_hd__dfrtp_4 _6349_ (.CLK(net91),
    .D(_0182_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[81] ));
 sky130_fd_sc_hd__dfrtp_2 _6350_ (.CLK(net92),
    .D(_0183_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[80] ));
 sky130_fd_sc_hd__dfxtp_1 _6351_ (.CLK(net93),
    .D(_0184_),
    .Q(\egd_top.BitStream_buffer.pc_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6352_ (.CLK(net94),
    .D(_0185_),
    .Q(\egd_top.BitStream_buffer.pc_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6353_ (.CLK(net95),
    .D(_0186_),
    .Q(\egd_top.BitStream_buffer.pc_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6354_ (.CLK(net96),
    .D(_0187_),
    .Q(\egd_top.BitStream_buffer.pc_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6355_ (.CLK(net97),
    .D(_0188_),
    .Q(\egd_top.BitStream_buffer.pc_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6356_ (.CLK(net98),
    .D(_0189_),
    .Q(\egd_top.BitStream_buffer.pc_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6357_ (.CLK(net99),
    .D(_0190_),
    .Q(\egd_top.BitStream_buffer.pc_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6358_ (.CLK(net100),
    .D(_0191_),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.BS_buffer[111] ));
 sky130_fd_sc_hd__dfrtp_1 _6359_ (.CLK(net101),
    .D(_0192_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[110] ));
 sky130_fd_sc_hd__dfrtp_1 _6360_ (.CLK(net102),
    .D(_0193_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[109] ));
 sky130_fd_sc_hd__dfrtp_1 _6361_ (.CLK(net103),
    .D(_0194_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[108] ));
 sky130_fd_sc_hd__dfrtp_1 _6362_ (.CLK(net104),
    .D(_0195_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[107] ));
 sky130_fd_sc_hd__dfrtp_1 _6363_ (.CLK(net105),
    .D(_0196_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[106] ));
 sky130_fd_sc_hd__dfrtp_1 _6364_ (.CLK(net106),
    .D(_0197_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[105] ));
 sky130_fd_sc_hd__dfrtp_1 _6365_ (.CLK(net107),
    .D(_0198_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[104] ));
 sky130_fd_sc_hd__dfrtp_1 _6366_ (.CLK(net108),
    .D(_0199_),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.BS_buffer[103] ));
 sky130_fd_sc_hd__dfrtp_1 _6367_ (.CLK(net109),
    .D(_0200_),
    .RESET_B(net42),
    .Q(\egd_top.BitStream_buffer.BS_buffer[102] ));
 sky130_fd_sc_hd__dfrtp_1 _6368_ (.CLK(net110),
    .D(_0201_),
    .RESET_B(net42),
    .Q(\egd_top.BitStream_buffer.BS_buffer[101] ));
 sky130_fd_sc_hd__dfrtp_1 _6369_ (.CLK(net111),
    .D(_0202_),
    .RESET_B(net42),
    .Q(\egd_top.BitStream_buffer.BS_buffer[100] ));
 sky130_fd_sc_hd__dfrtp_1 _6370_ (.CLK(net112),
    .D(_0203_),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.BS_buffer[99] ));
 sky130_fd_sc_hd__dfrtp_1 _6371_ (.CLK(net113),
    .D(_0204_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[98] ));
 sky130_fd_sc_hd__dfrtp_1 _6372_ (.CLK(net114),
    .D(_0205_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[97] ));
 sky130_fd_sc_hd__dfrtp_1 _6373_ (.CLK(net115),
    .D(_0206_),
    .RESET_B(net41),
    .Q(\egd_top.BitStream_buffer.BS_buffer[96] ));
 sky130_fd_sc_hd__dfrtp_2 _6374_ (.CLK(net116),
    .D(_0207_),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.buffer_index[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6375_ (.CLK(net117),
    .D(_0208_),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.buffer_index[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6376_ (.CLK(net118),
    .D(_0209_),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.buffer_index[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6377_ (.CLK(net119),
    .D(_0210_),
    .RESET_B(net51),
    .Q(\egd_top.BitStream_buffer.BS_buffer[79] ));
 sky130_fd_sc_hd__dfrtp_4 _6378_ (.CLK(net120),
    .D(_0211_),
    .RESET_B(net51),
    .Q(\egd_top.BitStream_buffer.BS_buffer[78] ));
 sky130_fd_sc_hd__dfrtp_4 _6379_ (.CLK(net121),
    .D(_0212_),
    .RESET_B(net51),
    .Q(\egd_top.BitStream_buffer.BS_buffer[77] ));
 sky130_fd_sc_hd__dfrtp_4 _6380_ (.CLK(net122),
    .D(_0213_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[76] ));
 sky130_fd_sc_hd__dfrtp_4 _6381_ (.CLK(net123),
    .D(_0214_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[75] ));
 sky130_fd_sc_hd__dfrtp_4 _6382_ (.CLK(net124),
    .D(_0215_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[74] ));
 sky130_fd_sc_hd__dfrtp_4 _6383_ (.CLK(net125),
    .D(_0216_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[73] ));
 sky130_fd_sc_hd__dfrtp_4 _6384_ (.CLK(net126),
    .D(_0217_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[72] ));
 sky130_fd_sc_hd__dfrtp_4 _6385_ (.CLK(net127),
    .D(_0218_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[71] ));
 sky130_fd_sc_hd__dfrtp_2 _6386_ (.CLK(net128),
    .D(_0219_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[70] ));
 sky130_fd_sc_hd__dfrtp_2 _6387_ (.CLK(net129),
    .D(_0220_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[69] ));
 sky130_fd_sc_hd__dfrtp_2 _6388_ (.CLK(net130),
    .D(_0221_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[68] ));
 sky130_fd_sc_hd__dfrtp_1 _6389_ (.CLK(net131),
    .D(_0222_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[67] ));
 sky130_fd_sc_hd__dfrtp_1 _6390_ (.CLK(net132),
    .D(_0223_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[66] ));
 sky130_fd_sc_hd__dfrtp_1 _6391_ (.CLK(net133),
    .D(_0224_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[65] ));
 sky130_fd_sc_hd__dfrtp_1 _6392_ (.CLK(net134),
    .D(_0225_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[64] ));
 sky130_fd_sc_hd__dfrtp_1 _6393_ (.CLK(net135),
    .D(_0226_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[63] ));
 sky130_fd_sc_hd__dfrtp_1 _6394_ (.CLK(net136),
    .D(_0227_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[62] ));
 sky130_fd_sc_hd__dfrtp_1 _6395_ (.CLK(net137),
    .D(_0228_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[61] ));
 sky130_fd_sc_hd__dfrtp_1 _6396_ (.CLK(net138),
    .D(_0229_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[60] ));
 sky130_fd_sc_hd__dfrtp_1 _6397_ (.CLK(net139),
    .D(_0230_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[59] ));
 sky130_fd_sc_hd__dfrtp_1 _6398_ (.CLK(net140),
    .D(_0231_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[58] ));
 sky130_fd_sc_hd__dfrtp_4 _6399_ (.CLK(net141),
    .D(_0232_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[57] ));
 sky130_fd_sc_hd__dfrtp_4 _6400_ (.CLK(net142),
    .D(_0233_),
    .RESET_B(net52),
    .Q(\egd_top.BitStream_buffer.BS_buffer[56] ));
 sky130_fd_sc_hd__dfrtp_4 _6401_ (.CLK(net143),
    .D(_0234_),
    .RESET_B(net52),
    .Q(\egd_top.BitStream_buffer.BS_buffer[55] ));
 sky130_fd_sc_hd__dfrtp_4 _6402_ (.CLK(net144),
    .D(_0235_),
    .RESET_B(net52),
    .Q(\egd_top.BitStream_buffer.BS_buffer[54] ));
 sky130_fd_sc_hd__dfrtp_4 _6403_ (.CLK(net145),
    .D(_0236_),
    .RESET_B(net52),
    .Q(\egd_top.BitStream_buffer.BS_buffer[53] ));
 sky130_fd_sc_hd__dfrtp_1 _6404_ (.CLK(net146),
    .D(_0237_),
    .RESET_B(net52),
    .Q(\egd_top.BitStream_buffer.BS_buffer[52] ));
 sky130_fd_sc_hd__dfrtp_1 _6405_ (.CLK(net147),
    .D(_0238_),
    .RESET_B(net52),
    .Q(\egd_top.BitStream_buffer.BS_buffer[51] ));
 sky130_fd_sc_hd__dfrtp_1 _6406_ (.CLK(net148),
    .D(_0239_),
    .RESET_B(net52),
    .Q(\egd_top.BitStream_buffer.BS_buffer[50] ));
 sky130_fd_sc_hd__dfrtp_1 _6407_ (.CLK(net149),
    .D(_0240_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[49] ));
 sky130_fd_sc_hd__dfrtp_1 _6408_ (.CLK(net150),
    .D(_0241_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[48] ));
 sky130_fd_sc_hd__dfrtp_1 _6409_ (.CLK(net151),
    .D(_0242_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[47] ));
 sky130_fd_sc_hd__dfrtp_4 _6410_ (.CLK(net152),
    .D(_0243_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[46] ));
 sky130_fd_sc_hd__dfrtp_1 _6411_ (.CLK(net153),
    .D(_0244_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[45] ));
 sky130_fd_sc_hd__dfrtp_1 _6412_ (.CLK(net154),
    .D(_0245_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[44] ));
 sky130_fd_sc_hd__dfrtp_1 _6413_ (.CLK(net155),
    .D(_0246_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[43] ));
 sky130_fd_sc_hd__dfrtp_1 _6414_ (.CLK(net156),
    .D(_0247_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[42] ));
 sky130_fd_sc_hd__dfrtp_1 _6415_ (.CLK(net157),
    .D(_0248_),
    .RESET_B(net48),
    .Q(\egd_top.BitStream_buffer.BS_buffer[41] ));
 sky130_fd_sc_hd__dfrtp_1 _6416_ (.CLK(net158),
    .D(_0249_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[40] ));
 sky130_fd_sc_hd__dfrtp_1 _6417_ (.CLK(net159),
    .D(_0250_),
    .RESET_B(net50),
    .Q(\egd_top.BitStream_buffer.BS_buffer[39] ));
 sky130_fd_sc_hd__dfrtp_1 _6418_ (.CLK(net160),
    .D(_0251_),
    .RESET_B(net49),
    .Q(\egd_top.BitStream_buffer.BS_buffer[38] ));
 sky130_fd_sc_hd__dfrtp_1 _6419_ (.CLK(net161),
    .D(_0252_),
    .RESET_B(net47),
    .Q(\egd_top.BitStream_buffer.BS_buffer[37] ));
 sky130_fd_sc_hd__dfrtp_1 _6420_ (.CLK(net162),
    .D(_0253_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[36] ));
 sky130_fd_sc_hd__dfrtp_1 _6421_ (.CLK(net163),
    .D(_0254_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[35] ));
 sky130_fd_sc_hd__dfrtp_1 _6422_ (.CLK(net164),
    .D(_0255_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[34] ));
 sky130_fd_sc_hd__dfrtp_1 _6423_ (.CLK(net165),
    .D(_0256_),
    .RESET_B(net41),
    .Q(\egd_top.BitStream_buffer.BS_buffer[33] ));
 sky130_fd_sc_hd__dfrtp_1 _6424_ (.CLK(net166),
    .D(_0257_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[32] ));
 sky130_fd_sc_hd__dfrtp_1 _6425_ (.CLK(net167),
    .D(_0258_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6426_ (.CLK(net168),
    .D(_0259_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[30] ));
 sky130_fd_sc_hd__dfrtp_1 _6427_ (.CLK(net169),
    .D(_0260_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[29] ));
 sky130_fd_sc_hd__dfrtp_1 _6428_ (.CLK(net170),
    .D(_0261_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[28] ));
 sky130_fd_sc_hd__dfrtp_1 _6429_ (.CLK(net171),
    .D(_0262_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[27] ));
 sky130_fd_sc_hd__dfrtp_1 _6430_ (.CLK(net172),
    .D(_0263_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[26] ));
 sky130_fd_sc_hd__dfrtp_1 _6431_ (.CLK(net173),
    .D(_0264_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[25] ));
 sky130_fd_sc_hd__dfrtp_1 _6432_ (.CLK(net174),
    .D(_0265_),
    .RESET_B(net41),
    .Q(\egd_top.BitStream_buffer.BS_buffer[24] ));
 sky130_fd_sc_hd__dfrtp_1 _6433_ (.CLK(net175),
    .D(_0266_),
    .RESET_B(net41),
    .Q(\egd_top.BitStream_buffer.BS_buffer[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6434_ (.CLK(net176),
    .D(_0267_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6435_ (.CLK(net177),
    .D(_0268_),
    .RESET_B(net41),
    .Q(\egd_top.BitStream_buffer.BS_buffer[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6436_ (.CLK(net178),
    .D(_0269_),
    .RESET_B(net40),
    .Q(\egd_top.BitStream_buffer.BS_buffer[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6437_ (.CLK(net179),
    .D(_0270_),
    .RESET_B(net41),
    .Q(\egd_top.BitStream_buffer.BS_buffer[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6438_ (.CLK(net180),
    .D(_0271_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6439_ (.CLK(net181),
    .D(_0272_),
    .RESET_B(net39),
    .Q(\egd_top.BitStream_buffer.BS_buffer[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6440_ (.CLK(net182),
    .D(_0273_),
    .RESET_B(net41),
    .Q(\egd_top.BitStream_buffer.BS_buffer[16] ));
 sky130_fd_sc_hd__dfrtp_1 _6441_ (.CLK(net183),
    .D(_0274_),
    .RESET_B(net42),
    .Q(\egd_top.BitStream_buffer.BS_buffer[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6442_ (.CLK(net184),
    .D(_0275_),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.BS_buffer[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6443_ (.CLK(net185),
    .D(_0276_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6444_ (.CLK(net186),
    .D(_0277_),
    .RESET_B(net46),
    .Q(\egd_top.BitStream_buffer.BS_buffer[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6445_ (.CLK(net187),
    .D(_0278_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6446_ (.CLK(net188),
    .D(_0279_),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.BS_buffer[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6447_ (.CLK(net189),
    .D(_0280_),
    .RESET_B(net38),
    .Q(\egd_top.BitStream_buffer.BS_buffer[9] ));
 sky130_fd_sc_hd__dfrtp_2 _6448_ (.CLK(net190),
    .D(_0281_),
    .RESET_B(net42),
    .Q(\egd_top.BitStream_buffer.BS_buffer[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6449_ (.CLK(net191),
    .D(_0282_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6450_ (.CLK(net192),
    .D(_0283_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6451_ (.CLK(net193),
    .D(_0284_),
    .RESET_B(net38),
    .Q(\egd_top.BitStream_buffer.BS_buffer[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6452_ (.CLK(net194),
    .D(_0285_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6453_ (.CLK(net195),
    .D(_0286_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6454_ (.CLK(net196),
    .D(_0287_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6455_ (.CLK(net197),
    .D(_0288_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BS_buffer[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6456_ (.CLK(net198),
    .D(_0289_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BS_buffer[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6457_ (.CLK(net199),
    .D(_0290_),
    .RESET_B(net38),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6458_ (.CLK(net200),
    .D(_0291_),
    .RESET_B(net38),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6459_ (.CLK(net201),
    .D(_0292_),
    .RESET_B(net38),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6460_ (.CLK(net202),
    .D(_0293_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6461_ (.CLK(net203),
    .D(_0294_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6462_ (.CLK(net204),
    .D(_0295_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6463_ (.CLK(net205),
    .D(_0296_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6464_ (.CLK(net206),
    .D(_0297_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6465_ (.CLK(net207),
    .D(_0298_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6466_ (.CLK(net208),
    .D(_0299_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6467_ (.CLK(net209),
    .D(_0300_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[11] ));
 sky130_fd_sc_hd__dfrtp_2 _6468_ (.CLK(net210),
    .D(_0301_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6469_ (.CLK(net211),
    .D(_0302_),
    .RESET_B(net43),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6470_ (.CLK(net212),
    .D(_0303_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6471_ (.CLK(net213),
    .D(_0304_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_output[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6472_ (.CLK(net214),
    .D(_0305_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[127] ));
 sky130_fd_sc_hd__dfrtp_4 _6473_ (.CLK(net215),
    .D(_0306_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[126] ));
 sky130_fd_sc_hd__dfrtp_4 _6474_ (.CLK(net216),
    .D(_0307_),
    .RESET_B(net44),
    .Q(\egd_top.BitStream_buffer.BS_buffer[125] ));
 sky130_fd_sc_hd__dfrtp_4 _6475_ (.CLK(net217),
    .D(_0308_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[124] ));
 sky130_fd_sc_hd__dfrtp_2 _6476_ (.CLK(net218),
    .D(_0309_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[123] ));
 sky130_fd_sc_hd__dfrtp_2 _6477_ (.CLK(net219),
    .D(_0310_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[122] ));
 sky130_fd_sc_hd__dfrtp_1 _6478_ (.CLK(net220),
    .D(_0311_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[121] ));
 sky130_fd_sc_hd__dfrtp_1 _6479_ (.CLK(net53),
    .D(_0312_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[120] ));
 sky130_fd_sc_hd__dfrtp_1 _6480_ (.CLK(net54),
    .D(_0313_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[119] ));
 sky130_fd_sc_hd__dfrtp_1 _6481_ (.CLK(net55),
    .D(_0314_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[118] ));
 sky130_fd_sc_hd__dfrtp_1 _6482_ (.CLK(net56),
    .D(_0315_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[117] ));
 sky130_fd_sc_hd__dfrtp_1 _6483_ (.CLK(net57),
    .D(_0316_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[116] ));
 sky130_fd_sc_hd__dfrtp_1 _6484_ (.CLK(net58),
    .D(_0317_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[115] ));
 sky130_fd_sc_hd__dfrtp_1 _6485_ (.CLK(net59),
    .D(_0318_),
    .RESET_B(net45),
    .Q(\egd_top.BitStream_buffer.BS_buffer[114] ));
 sky130_fd_sc_hd__dfrtp_1 _6486_ (.CLK(net60),
    .D(_0319_),
    .RESET_B(net46),
    .Q(\egd_top.BitStream_buffer.BS_buffer[113] ));
 sky130_fd_sc_hd__dfrtp_1 _6487_ (.CLK(net61),
    .D(_0320_),
    .RESET_B(net46),
    .Q(\egd_top.BitStream_buffer.BS_buffer[112] ));
 sky130_fd_sc_hd__dfstp_1 _6488_ (.CLK(net62),
    .D(_0321_),
    .SET_B(net38),
    .Q(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ));
 sky130_fd_sc_hd__dfrtp_4 _6489_ (.CLK(net63),
    .D(_0322_),
    .RESET_B(net36),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_4 _6490_ (.CLK(net64),
    .D(_0323_),
    .RESET_B(net36),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_4 _6491_ (.CLK(net65),
    .D(_0324_),
    .RESET_B(net35),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _6492_ (.CLK(net66),
    .D(\egd_top.BitStream_buffer.pc[0] ),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.pc_previous[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6493_ (.CLK(net67),
    .D(\egd_top.BitStream_buffer.pc[1] ),
    .RESET_B(net37),
    .Q(\egd_top.BitStream_buffer.pc_previous[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6494_ (.CLK(net68),
    .D(\egd_top.BitStream_buffer.pc[2] ),
    .RESET_B(net36),
    .Q(\egd_top.BitStream_buffer.pc_previous[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6495_ (.CLK(net69),
    .D(\egd_top.BitStream_buffer.pc[3] ),
    .RESET_B(net36),
    .Q(\egd_top.BitStream_buffer.pc_previous[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6496_ (.CLK(net70),
    .D(\egd_top.BitStream_buffer.pc[4] ),
    .RESET_B(net36),
    .Q(\egd_top.BitStream_buffer.pc_previous[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6497_ (.CLK(net71),
    .D(\egd_top.BitStream_buffer.pc[5] ),
    .RESET_B(net36),
    .Q(\egd_top.BitStream_buffer.pc_previous[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6498_ (.CLK(net72),
    .D(\egd_top.BitStream_buffer.pc[6] ),
    .RESET_B(net35),
    .Q(\egd_top.BitStream_buffer.pc_previous[6] ));
 sky130_fd_sc_hd__dfrtp_2 _6499_ (.CLK(net73),
    .D(_0325_),
    .RESET_B(net35),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_4 _6500_ (.CLK(net74),
    .D(_0326_),
    .RESET_B(net39),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_2 _6501_ (.CLK(net75),
    .D(_0327_),
    .RESET_B(net39),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_2 _6502_ (.CLK(net76),
    .D(_0328_),
    .RESET_B(net39),
    .Q(net34));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2717_ (.A(_2717_),
    .X(clknet_0__2717_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2718_ (.A(_2718_),
    .X(clknet_0__2718_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2719_ (.A(_2719_),
    .X(clknet_0__2719_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2720_ (.A(_2720_),
    .X(clknet_0__2720_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2721_ (.A(_2721_),
    .X(clknet_0__2721_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2722_ (.A(_2722_),
    .X(clknet_0__2722_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2723_ (.A(_2723_),
    .X(clknet_0__2723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2724_ (.A(_2724_),
    .X(clknet_0__2724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2725_ (.A(_2725_),
    .X(clknet_0__2725_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2726_ (.A(_2726_),
    .X(clknet_0__2726_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2727_ (.A(_2727_),
    .X(clknet_0__2727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2728_ (.A(_2728_),
    .X(clknet_0__2728_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2729_ (.A(_2729_),
    .X(clknet_0__2729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2730_ (.A(_2730_),
    .X(clknet_0__2730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__2731_ (.A(_2731_),
    .X(clknet_0__2731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2717_ (.A(clknet_0__2717_),
    .X(clknet_1_0__leaf__2717_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2718_ (.A(clknet_0__2718_),
    .X(clknet_1_0__leaf__2718_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2719_ (.A(clknet_0__2719_),
    .X(clknet_1_0__leaf__2719_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2720_ (.A(clknet_0__2720_),
    .X(clknet_1_0__leaf__2720_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2721_ (.A(clknet_0__2721_),
    .X(clknet_1_0__leaf__2721_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2722_ (.A(clknet_0__2722_),
    .X(clknet_1_0__leaf__2722_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2723_ (.A(clknet_0__2723_),
    .X(clknet_1_0__leaf__2723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2724_ (.A(clknet_0__2724_),
    .X(clknet_1_0__leaf__2724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2725_ (.A(clknet_0__2725_),
    .X(clknet_1_0__leaf__2725_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2726_ (.A(clknet_0__2726_),
    .X(clknet_1_0__leaf__2726_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2727_ (.A(clknet_0__2727_),
    .X(clknet_1_0__leaf__2727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2728_ (.A(clknet_0__2728_),
    .X(clknet_1_0__leaf__2728_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2729_ (.A(clknet_0__2729_),
    .X(clknet_1_0__leaf__2729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2730_ (.A(clknet_0__2730_),
    .X(clknet_1_0__leaf__2730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__2731_ (.A(clknet_0__2731_),
    .X(clknet_1_0__leaf__2731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2717_ (.A(clknet_0__2717_),
    .X(clknet_1_1__leaf__2717_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2718_ (.A(clknet_0__2718_),
    .X(clknet_1_1__leaf__2718_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2719_ (.A(clknet_0__2719_),
    .X(clknet_1_1__leaf__2719_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2720_ (.A(clknet_0__2720_),
    .X(clknet_1_1__leaf__2720_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2721_ (.A(clknet_0__2721_),
    .X(clknet_1_1__leaf__2721_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2722_ (.A(clknet_0__2722_),
    .X(clknet_1_1__leaf__2722_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2723_ (.A(clknet_0__2723_),
    .X(clknet_1_1__leaf__2723_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2724_ (.A(clknet_0__2724_),
    .X(clknet_1_1__leaf__2724_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2725_ (.A(clknet_0__2725_),
    .X(clknet_1_1__leaf__2725_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2726_ (.A(clknet_0__2726_),
    .X(clknet_1_1__leaf__2726_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2727_ (.A(clknet_0__2727_),
    .X(clknet_1_1__leaf__2727_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2728_ (.A(clknet_0__2728_),
    .X(clknet_1_1__leaf__2728_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2729_ (.A(clknet_0__2729_),
    .X(clknet_1_1__leaf__2729_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2730_ (.A(clknet_0__2730_),
    .X(clknet_1_1__leaf__2730_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__2731_ (.A(clknet_0__2731_),
    .X(clknet_1_1__leaf__2731_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__buf_4 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net46),
    .X(net36));
 sky130_fd_sc_hd__buf_4 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net46),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net41),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net46),
    .X(net42));
 sky130_fd_sc_hd__buf_4 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net19),
    .X(net46));
 sky130_fd_sc_hd__buf_4 fanout47 (.A(net51),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__buf_4 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_2 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net19),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1 (.A(net225),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net34),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_2792_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_2793_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\egd_top.BitStream_buffer.BitStream_buffer_valid_n ),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(la_data_in_47_32[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(la_data_in_47_32[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(la_data_in_47_32[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(la_data_in_47_32[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(la_data_in_47_32[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(la_data_in_47_32[7]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(la_data_in_47_32[8]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(la_data_in_47_32[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(la_data_in_49_48[0]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(la_data_in_49_48[1]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(la_data_in_65),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(la_data_in_47_32[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input3 (.A(la_data_in_47_32[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(la_data_in_47_32[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(la_data_in_47_32[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(la_data_in_47_32[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(la_data_in_47_32[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(la_data_in_47_32[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(la_data_in_47_32[2]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(la_data_out_15_8[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(la_data_out_15_8[1]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(la_data_out_15_8[2]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(la_data_out_15_8[3]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(la_data_out_15_8[4]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(la_data_out_15_8[5]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(la_data_out_15_8[6]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(la_data_out_15_8[7]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(la_data_out_18_16[0]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(la_data_out_18_16[1]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(la_data_out_18_16[2]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(la_data_out_22_19[0]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(la_data_out_22_19[1]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(la_data_out_22_19[2]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(la_data_out_22_19[3]));
endmodule

