magic
tech sky130A
magscale 1 2
timestamp 1697107604
<< obsli1 >>
rect 1104 2159 52348 53329
<< obsm1 >>
rect 934 1980 53162 53360
<< metal2 >>
rect 1674 0 1730 800
rect 3238 0 3294 800
rect 4802 0 4858 800
rect 6366 0 6422 800
rect 7930 0 7986 800
rect 9494 0 9550 800
rect 11058 0 11114 800
rect 12622 0 12678 800
rect 14186 0 14242 800
rect 15750 0 15806 800
rect 17314 0 17370 800
rect 18878 0 18934 800
rect 20442 0 20498 800
rect 22006 0 22062 800
rect 23570 0 23626 800
rect 25134 0 25190 800
rect 26698 0 26754 800
rect 28262 0 28318 800
rect 29826 0 29882 800
rect 31390 0 31446 800
rect 32954 0 33010 800
rect 34518 0 34574 800
rect 36082 0 36138 800
rect 37646 0 37702 800
rect 39210 0 39266 800
rect 40774 0 40830 800
rect 42338 0 42394 800
rect 43902 0 43958 800
rect 45466 0 45522 800
rect 47030 0 47086 800
rect 48594 0 48650 800
rect 50158 0 50214 800
rect 51722 0 51778 800
<< obsm2 >>
rect 938 856 53156 53349
rect 938 734 1618 856
rect 1786 734 3182 856
rect 3350 734 4746 856
rect 4914 734 6310 856
rect 6478 734 7874 856
rect 8042 734 9438 856
rect 9606 734 11002 856
rect 11170 734 12566 856
rect 12734 734 14130 856
rect 14298 734 15694 856
rect 15862 734 17258 856
rect 17426 734 18822 856
rect 18990 734 20386 856
rect 20554 734 21950 856
rect 22118 734 23514 856
rect 23682 734 25078 856
rect 25246 734 26642 856
rect 26810 734 28206 856
rect 28374 734 29770 856
rect 29938 734 31334 856
rect 31502 734 32898 856
rect 33066 734 34462 856
rect 34630 734 36026 856
rect 36194 734 37590 856
rect 37758 734 39154 856
rect 39322 734 40718 856
rect 40886 734 42282 856
rect 42450 734 43846 856
rect 44014 734 45410 856
rect 45578 734 46974 856
rect 47142 734 48538 856
rect 48706 734 50102 856
rect 50270 734 51666 856
rect 51834 734 53156 856
<< metal3 >>
rect 0 41624 800 41744
rect 0 13880 800 14000
<< obsm3 >>
rect 800 41824 52887 53345
rect 880 41544 52887 41824
rect 800 14080 52887 41544
rect 880 13800 52887 14080
rect 800 2143 52887 13800
<< metal4 >>
rect 4208 2128 4528 53360
rect 19568 2128 19888 53360
rect 34928 2128 35248 53360
rect 50288 2128 50608 53360
<< obsm4 >>
rect 6499 3435 19488 48653
rect 19968 3435 34848 48653
rect 35328 3435 50208 48653
rect 50688 3435 50909 48653
<< labels >>
rlabel metal2 s 25134 0 25190 800 6 la_data_in_47_32[0]
port 1 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in_47_32[10]
port 2 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in_47_32[11]
port 3 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in_47_32[12]
port 4 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in_47_32[13]
port 5 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in_47_32[14]
port 6 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in_47_32[15]
port 7 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_data_in_47_32[1]
port 8 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in_47_32[2]
port 9 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 la_data_in_47_32[3]
port 10 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in_47_32[4]
port 11 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_data_in_47_32[5]
port 12 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in_47_32[6]
port 13 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in_47_32[7]
port 14 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_data_in_47_32[8]
port 15 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in_47_32[9]
port 16 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_data_in_49_48[0]
port 17 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_data_in_49_48[1]
port 18 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 la_data_out_15_8[0]
port 19 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 la_data_out_15_8[1]
port 20 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 la_data_out_15_8[2]
port 21 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 la_data_out_15_8[3]
port 22 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 la_data_out_15_8[4]
port 23 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 la_data_out_15_8[5]
port 24 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 la_data_out_15_8[6]
port 25 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 la_data_out_15_8[7]
port 26 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 la_data_out_18_16[0]
port 27 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 la_data_out_18_16[1]
port 28 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 la_data_out_18_16[2]
port 29 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 la_data_out_22_19[0]
port 30 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 la_data_out_22_19[1]
port 31 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 la_data_out_22_19[2]
port 32 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 la_data_out_22_19[3]
port 33 nsew signal output
rlabel metal4 s 4208 2128 4528 53360 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 53360 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 53360 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 53360 6 vssd1
port 35 nsew ground bidirectional
rlabel metal3 s 0 13880 800 14000 6 wb_clk_i
port 36 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 wb_rst_i
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 53460 55604
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10109206
string GDS_FILE /home/uniccass/H.264_Decoder/openlane/egd_top_wrapper/runs/23_10_12_03_22/results/signoff/egd_top_wrapper.magic.gds
string GDS_START 676554
<< end >>

