VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO egd_top
  CLASS BLOCK ;
  FOREIGN egd_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 249.865 BY 260.585 ;
  PIN BitStream_buffer_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END BitStream_buffer_input[0]
  PIN BitStream_buffer_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END BitStream_buffer_input[10]
  PIN BitStream_buffer_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END BitStream_buffer_input[11]
  PIN BitStream_buffer_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END BitStream_buffer_input[12]
  PIN BitStream_buffer_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END BitStream_buffer_input[13]
  PIN BitStream_buffer_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END BitStream_buffer_input[14]
  PIN BitStream_buffer_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END BitStream_buffer_input[15]
  PIN BitStream_buffer_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END BitStream_buffer_input[1]
  PIN BitStream_buffer_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END BitStream_buffer_input[2]
  PIN BitStream_buffer_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END BitStream_buffer_input[3]
  PIN BitStream_buffer_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END BitStream_buffer_input[4]
  PIN BitStream_buffer_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END BitStream_buffer_input[5]
  PIN BitStream_buffer_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END BitStream_buffer_input[6]
  PIN BitStream_buffer_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END BitStream_buffer_input[7]
  PIN BitStream_buffer_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END BitStream_buffer_input[8]
  PIN BitStream_buffer_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END BitStream_buffer_input[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END clk
  PIN exp_golomb_decoding_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END exp_golomb_decoding_output[0]
  PIN exp_golomb_decoding_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END exp_golomb_decoding_output[1]
  PIN exp_golomb_decoding_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END exp_golomb_decoding_output[2]
  PIN exp_golomb_decoding_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END exp_golomb_decoding_output[3]
  PIN exp_golomb_decoding_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END exp_golomb_decoding_output[4]
  PIN exp_golomb_decoding_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END exp_golomb_decoding_output[5]
  PIN exp_golomb_decoding_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END exp_golomb_decoding_output[6]
  PIN exp_golomb_decoding_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END exp_golomb_decoding_output[7]
  PIN exp_golomb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END exp_golomb_sel[0]
  PIN exp_golomb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END exp_golomb_sel[1]
  PIN half_fill_counter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END half_fill_counter[0]
  PIN half_fill_counter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END half_fill_counter[1]
  PIN half_fill_counter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END half_fill_counter[2]
  PIN reset_counter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END reset_counter[0]
  PIN reset_counter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END reset_counter[1]
  PIN reset_counter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END reset_counter[2]
  PIN reset_counter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END reset_counter[3]
  PIN reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END reset_n
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 247.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 247.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 247.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 246.105 244.450 247.710 ;
        RECT 5.330 240.665 244.450 243.495 ;
        RECT 5.330 235.225 244.450 238.055 ;
        RECT 5.330 229.785 244.450 232.615 ;
        RECT 5.330 224.345 244.450 227.175 ;
        RECT 5.330 218.905 244.450 221.735 ;
        RECT 5.330 213.465 244.450 216.295 ;
        RECT 5.330 208.025 244.450 210.855 ;
        RECT 5.330 202.585 244.450 205.415 ;
        RECT 5.330 197.145 244.450 199.975 ;
        RECT 5.330 191.705 244.450 194.535 ;
        RECT 5.330 186.265 244.450 189.095 ;
        RECT 5.330 180.825 244.450 183.655 ;
        RECT 5.330 175.385 244.450 178.215 ;
        RECT 5.330 169.945 244.450 172.775 ;
        RECT 5.330 164.505 244.450 167.335 ;
        RECT 5.330 159.065 244.450 161.895 ;
        RECT 5.330 153.625 244.450 156.455 ;
        RECT 5.330 148.185 244.450 151.015 ;
        RECT 5.330 142.745 244.450 145.575 ;
        RECT 5.330 137.305 244.450 140.135 ;
        RECT 5.330 131.865 244.450 134.695 ;
        RECT 5.330 126.425 244.450 129.255 ;
        RECT 5.330 120.985 244.450 123.815 ;
        RECT 5.330 115.545 244.450 118.375 ;
        RECT 5.330 110.105 244.450 112.935 ;
        RECT 5.330 104.665 244.450 107.495 ;
        RECT 5.330 99.225 244.450 102.055 ;
        RECT 5.330 93.785 244.450 96.615 ;
        RECT 5.330 88.345 244.450 91.175 ;
        RECT 5.330 82.905 244.450 85.735 ;
        RECT 5.330 77.465 244.450 80.295 ;
        RECT 5.330 72.025 244.450 74.855 ;
        RECT 5.330 66.585 244.450 69.415 ;
        RECT 5.330 61.145 244.450 63.975 ;
        RECT 5.330 55.705 244.450 58.535 ;
        RECT 5.330 50.265 244.450 53.095 ;
        RECT 5.330 44.825 244.450 47.655 ;
        RECT 5.330 39.385 244.450 42.215 ;
        RECT 5.330 33.945 244.450 36.775 ;
        RECT 5.330 28.505 244.450 31.335 ;
        RECT 5.330 23.065 244.450 25.895 ;
        RECT 5.330 17.625 244.450 20.455 ;
        RECT 5.330 12.185 244.450 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 244.260 247.605 ;
      LAYER met1 ;
        RECT 5.520 7.520 244.260 247.760 ;
      LAYER met2 ;
        RECT 7.000 4.280 242.260 247.705 ;
        RECT 7.000 3.670 7.170 4.280 ;
        RECT 8.010 3.670 14.070 4.280 ;
        RECT 14.910 3.670 20.970 4.280 ;
        RECT 21.810 3.670 27.870 4.280 ;
        RECT 28.710 3.670 34.770 4.280 ;
        RECT 35.610 3.670 41.670 4.280 ;
        RECT 42.510 3.670 48.570 4.280 ;
        RECT 49.410 3.670 55.470 4.280 ;
        RECT 56.310 3.670 62.370 4.280 ;
        RECT 63.210 3.670 69.270 4.280 ;
        RECT 70.110 3.670 76.170 4.280 ;
        RECT 77.010 3.670 83.070 4.280 ;
        RECT 83.910 3.670 89.970 4.280 ;
        RECT 90.810 3.670 96.870 4.280 ;
        RECT 97.710 3.670 103.770 4.280 ;
        RECT 104.610 3.670 110.670 4.280 ;
        RECT 111.510 3.670 117.570 4.280 ;
        RECT 118.410 3.670 124.470 4.280 ;
        RECT 125.310 3.670 131.370 4.280 ;
        RECT 132.210 3.670 138.270 4.280 ;
        RECT 139.110 3.670 145.170 4.280 ;
        RECT 146.010 3.670 152.070 4.280 ;
        RECT 152.910 3.670 158.970 4.280 ;
        RECT 159.810 3.670 165.870 4.280 ;
        RECT 166.710 3.670 172.770 4.280 ;
        RECT 173.610 3.670 179.670 4.280 ;
        RECT 180.510 3.670 186.570 4.280 ;
        RECT 187.410 3.670 193.470 4.280 ;
        RECT 194.310 3.670 200.370 4.280 ;
        RECT 201.210 3.670 207.270 4.280 ;
        RECT 208.110 3.670 214.170 4.280 ;
        RECT 215.010 3.670 221.070 4.280 ;
        RECT 221.910 3.670 227.970 4.280 ;
        RECT 228.810 3.670 234.870 4.280 ;
        RECT 235.710 3.670 241.770 4.280 ;
      LAYER met3 ;
        RECT 12.485 8.350 241.895 247.685 ;
      LAYER met4 ;
        RECT 16.855 11.055 20.640 173.225 ;
        RECT 23.040 11.055 97.440 173.225 ;
        RECT 99.840 11.055 174.240 173.225 ;
        RECT 176.640 11.055 220.505 173.225 ;
  END
END egd_top
END LIBRARY

