VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO egd_top_wrapper
  CLASS BLOCK ;
  FOREIGN egd_top_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 259.975 BY 270.695 ;
  PIN la_data_in_47_32[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END la_data_in_47_32[0]
  PIN la_data_in_47_32[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END la_data_in_47_32[10]
  PIN la_data_in_47_32[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END la_data_in_47_32[11]
  PIN la_data_in_47_32[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END la_data_in_47_32[12]
  PIN la_data_in_47_32[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END la_data_in_47_32[13]
  PIN la_data_in_47_32[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END la_data_in_47_32[14]
  PIN la_data_in_47_32[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END la_data_in_47_32[15]
  PIN la_data_in_47_32[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END la_data_in_47_32[1]
  PIN la_data_in_47_32[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END la_data_in_47_32[2]
  PIN la_data_in_47_32[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END la_data_in_47_32[3]
  PIN la_data_in_47_32[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END la_data_in_47_32[4]
  PIN la_data_in_47_32[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END la_data_in_47_32[5]
  PIN la_data_in_47_32[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END la_data_in_47_32[6]
  PIN la_data_in_47_32[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END la_data_in_47_32[7]
  PIN la_data_in_47_32[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END la_data_in_47_32[8]
  PIN la_data_in_47_32[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END la_data_in_47_32[9]
  PIN la_data_in_49_48[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END la_data_in_49_48[0]
  PIN la_data_in_49_48[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END la_data_in_49_48[1]
  PIN la_data_in_64
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_data_in_64
  PIN la_data_in_65
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_in_65
  PIN la_data_out_15_8[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END la_data_out_15_8[0]
  PIN la_data_out_15_8[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END la_data_out_15_8[1]
  PIN la_data_out_15_8[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END la_data_out_15_8[2]
  PIN la_data_out_15_8[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END la_data_out_15_8[3]
  PIN la_data_out_15_8[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END la_data_out_15_8[4]
  PIN la_data_out_15_8[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END la_data_out_15_8[5]
  PIN la_data_out_15_8[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END la_data_out_15_8[6]
  PIN la_data_out_15_8[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END la_data_out_15_8[7]
  PIN la_data_out_18_16[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END la_data_out_18_16[0]
  PIN la_data_out_18_16[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END la_data_out_18_16[1]
  PIN la_data_out_18_16[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END la_data_out_18_16[2]
  PIN la_data_out_22_19[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END la_data_out_22_19[0]
  PIN la_data_out_22_19[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END la_data_out_22_19[1]
  PIN la_data_out_22_19[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END la_data_out_22_19[2]
  PIN la_data_out_22_19[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END la_data_out_22_19[3]
  PIN la_oenb_64
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END la_oenb_64
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 258.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 258.640 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 258.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 258.640 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 254.380 258.485 ;
      LAYER met1 ;
        RECT 5.520 6.840 254.380 258.640 ;
      LAYER met2 ;
        RECT 8.840 4.280 254.280 258.585 ;
        RECT 9.390 3.670 15.450 4.280 ;
        RECT 16.290 3.670 22.350 4.280 ;
        RECT 23.190 3.670 29.250 4.280 ;
        RECT 30.090 3.670 36.150 4.280 ;
        RECT 36.990 3.670 43.050 4.280 ;
        RECT 43.890 3.670 49.950 4.280 ;
        RECT 50.790 3.670 56.850 4.280 ;
        RECT 57.690 3.670 63.750 4.280 ;
        RECT 64.590 3.670 70.650 4.280 ;
        RECT 71.490 3.670 77.550 4.280 ;
        RECT 78.390 3.670 84.450 4.280 ;
        RECT 85.290 3.670 91.350 4.280 ;
        RECT 92.190 3.670 98.250 4.280 ;
        RECT 99.090 3.670 105.150 4.280 ;
        RECT 105.990 3.670 112.050 4.280 ;
        RECT 112.890 3.670 118.950 4.280 ;
        RECT 119.790 3.670 125.850 4.280 ;
        RECT 126.690 3.670 132.750 4.280 ;
        RECT 133.590 3.670 139.650 4.280 ;
        RECT 140.490 3.670 146.550 4.280 ;
        RECT 147.390 3.670 153.450 4.280 ;
        RECT 154.290 3.670 160.350 4.280 ;
        RECT 161.190 3.670 167.250 4.280 ;
        RECT 168.090 3.670 174.150 4.280 ;
        RECT 174.990 3.670 181.050 4.280 ;
        RECT 181.890 3.670 187.950 4.280 ;
        RECT 188.790 3.670 194.850 4.280 ;
        RECT 195.690 3.670 201.750 4.280 ;
        RECT 202.590 3.670 208.650 4.280 ;
        RECT 209.490 3.670 215.550 4.280 ;
        RECT 216.390 3.670 222.450 4.280 ;
        RECT 223.290 3.670 229.350 4.280 ;
        RECT 230.190 3.670 236.250 4.280 ;
        RECT 237.090 3.670 243.150 4.280 ;
        RECT 243.990 3.670 250.050 4.280 ;
        RECT 250.890 3.670 254.280 4.280 ;
      LAYER met3 ;
        RECT 4.000 135.680 253.855 258.565 ;
        RECT 4.400 134.280 253.855 135.680 ;
        RECT 4.000 9.695 253.855 134.280 ;
      LAYER met4 ;
        RECT 46.295 10.375 97.440 221.505 ;
        RECT 99.840 10.375 174.240 221.505 ;
        RECT 176.640 10.375 244.425 221.505 ;
  END
END egd_top_wrapper
END LIBRARY

